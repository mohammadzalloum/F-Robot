PK   e*X���H&  C�    cirkitFile.json�}ے�6r��(J�fq"ȹ��v��w�X9�3<J��=��^����e�LN�]<��X�����\H�MH"�<|@��������M���z�~~Z��n�c��~�O�߭>����?l��?����~��?��������i�7i)�TFy.m�c�Gy�%Q\d2�mZԕx�W���;�u�{]�^W��5�>�rш�溊���E�F�*��4u)UY�v_��pF�9#'���4yel�����D�Jd$�5�,u�Mcd�YJ��)kh�:c͚p��6��%kl���۷�����zݯN1�y�+ϼeF7q-Md�:�tm���?U�i[VFV��#�41��F�6����(��2�%џ%��
�jk��Z�F�M�&M�*��RՑ�RFER4�nd&�>IHb��*/u��}�0�V&�w�<"b
]Թ�4[�wS�c���&�"-h'HuZF�&j��*�pb��nLeS	�ѸR�Qj�4�!E,k)L�{7!����H��*�}�(��(Mem�I�U�P�M3dlA4�:ҙ)�4�27����kߖ	�d��]H@<�BK�#Ԑp�py�-�Dm�HĖޭ�:���D2n�<���Ļ�􌛖u뜦I�؍K��41�ʴHӆ�H}�Ʀ�Y]�IuB�\Q��"2R��q�$�b-�I��-�9	���FΘۣϢ�u��$^�M
bWE;Fj�**ˢ��F�{����&��Q��mZFQ�(A&����$�~����߾	���Ɔ�Lҙ�_$��}N�QÆ��RD%��[�sZ�]�5���p�����[�����/��5gh�z ]k��,�?c����5gl�E
Y<9�)4hh���)4�.�}�O�A. kh�Sh�%��`C��4���w>�����=��H���$��q�]�Q�����c]���H�֊^�+��U$&M�,6�I��+����X2c��8�d~6R��U��2�2ˣ2U&3�J��}����<c�<�)0fs�6�	8�E�~�!C'��s����i��"�[IMr�G�4	h.��mbx�� 24�o���}�C{10ft>C#�C�`\�A�ϊ9=>2(c��}6$���G�~f����7׼�|�Q�[����@���?�!��n�[���ڷ@��}K��˂^�����9s����j�=��#л�V��ڧ� �ٷ:�<��04�o]B^�oY��(a�lF��7۠[y�2��] �.�l��C�-�k"0z�P�s�@���Q�D��^!�s��"*K��Ma���EdS�,7yY뉘����&�fdW�Add�pC.�����@�l�����4\@ �}��Ti���n�jȩU5�69m�������T�_���&��i�TqEdǍ��������w�z��)�iv���}84��rh����l��Ai�-���~Kfq�"�Y��}."��f 10��S�����.0g���04������'B���loLK�\��Q���c���<��1F��-�o5�EB� "����������V����a�Z}��<@V�W�^d�^T�^��iȟ���-��F/��%��F/�������K��"Ө��K����� |>���u�{��Q#�F�q����h��8N="� �_�P�^f$z*�1��ܓ]@O�L/�$H�/Jv�ت�@�lZ����2��da�n/�6iN7���&�xԄ_����dAM	I�n��Cէ�v>�9�� �a�)��m�bntNI3�s�8��׵!uÚ�V���Rg�����X��t[)N�T&%g�m�8KҼN9��8m�a8���(�u�(G�Ӗ
���ʜ�$P���%�}�%W_�2-3��"�gE1N��H���P`ⴅ��̮��4
���8�i�7�i���Y�	���E��]@7�	�X�iŵ�;G
7��E�Mo�(��Y��iB�`ӫv��֩��BAZӫ\Mӂ���-5my���iN� �i�EqJ�� 
9��>4-�(h��%>�����v@��4-(���n���:3�P�4-(�ezvQx��E�{V#5�^G(�d�x2�B1$Ӵ�P� ���E��$s@��t� �{LG	P���
@aӁVQ1c����/BA�1kYU�s���{�r����#��� � ����h�?@/��'��?�z߲�/�|[s��O��v�?2���^d�^T�^t�^L�^� �� ��Az��H] �#wbv�Yu~/ah��8���evA�Yu~/�Ϊ�{�]�pV=���0�;���z�n��#�"��02,��#�2��@:8��0R,�H�#�2��0R,�H�#�*��Y)����^fi����^��2���:���/����^f�Ϊ�{�՜pV��ˬބ���^f9g�'{����^f�Ϊ�{��:8���eV��:��ٽΪ�{��8���eV^�:��Yy����^fyg��� ��U����Yم���^feΪO��hV���,��:��YZ�:���5�f�����g�����g���̧�Ь:��0�̧	Ь�d/pV��˼��f������hV��KZ�}X4���e��D���;,�U��2o��Y�C/��я��N�?����ޙ��O�M�����6��a�������{V�Vp���t+���u�Ȱ�f�$��9���d���<C��Z��3�޲n��k���X�4�G{
C�7�p��D�=#s����pʤ��;���P?'x����p���"�#8#{������.X��G���5�g�g�3߷�f���ɓ�+0��L@q�J�����v����9��X0�Мe�.���t"����1��[�%f�<#s�)���0��32���d�.�j�1�=V7\C"�K	��. a`>��̪yg��py��}�zQ~pS�>Fc�>Nj��.ɹf�����S�,�w��C�e�9��s��Rc��؁YG��^/=A��-�i,wv�}�'��l��aI5�t�~�"��f7�2��.����`⟣LX9Cn��z̿�/�L�*Գ[�T(K{�6j�����/��`X �:�0 !�G�/.�^���siy�� �XC{�  �XC{o%���ڗWa}�U������?=����j�󞈼!$��G��.@�O�ç�י��*��I
���3����� �ß&��/�L`�$����	��|&)�ڇO �s1)D�?|��I���O�Rp�����)������F�p
���F�b� �j]L���I�ܚ$�����¸�p�\|
����-D��GcB�.�
P��$� |1��� �+Ȏ��Mp����d��B&�b��v1!D�iSD(Dm�W@��)`�.&�(nmZ� _��&BQl��5>f7���b���S0�u�8w�6	�7I�5�~L&H�~,ū�����D&q:\t$���  �r�k����x9D)^�4C������E\��D��*j`*}pe<�']�y[}|ܓF����bF�c�]�@�/_�z��	�r�\��N�J����P'�j���P~�U�7�T&u�U҉|1��rA(r���C�r1��+X��P��*�� 0�_�R���~)}�w>j��ǻU��^�O�
��ߟuX]���u�-���
�����b��nU���|�6Z-�םm���u�Y\p��^w�$<\H�ם��2ZQ�ם��1\Z����֢�����u�Q+S;��'V2��O���SF6�\�a~��J���Lr�K��͸�7\���Y[�;\�#���@�%�+�m�IV#��GC��L3l��d��~�:�x��#�Gˡ����l j��Q� ���sLׇb�ˈ�g��p}�N������S��!<���Nw#���pE�^w�¥11��52{�y��Xf�:|����Σ��+�:����5=�6\J�7Y-��8�C���ʦg�����(��61Q�+n�n��nr��L�I���Y�L�uW��L�и��������9�3\(�s�bĒ�P7"Y�u��Ė1\��.�٣γ*�*���<�.�	
\�ӳ���=r8I�����ŗ\��������up�^w�	.��*�2(F\"c\+�G�g����z)\.��>\(��9��C=���B9��܁˅�zh��9��P���0p�Ple�5D{�	���D}VZF�:��h��8 �)�-)�#��G7g��h�;cds��=�9��Gv���pE�noB�Ҥoݬ+ݠ�_vI�޽_9��$��!n{vKݩZ'6nq4�ihCumŁ��.]޿8�ڶ٬օl����n]��yh��v��FTk\����*Z���
Z�e��A+$��F�G��|H���lD
;� �(��aF�άRH�g@&����:B\KGw罿΄!Y���$��;#"�r煲)�B4}��;v�lT�պ��-��Z�nw� [��b-v^@̻���3d��X������]hRV��[���_w����:E��cuo+i���:b����9���Ô+�v=�aF�A�D�0_Π�]�z���*W��I8s���$'�ˉ�q���Z�z\|0$�BqR����pS�����$����9`NN���8�C��|�Ŏ8 N֙��s��-'�Ɖ�q���'Z�	��\��ݫ\�=��g�^���1>c�y��W)�>0lK1W��=Ĉ��u�|0jؕ�����-�=D5�Ss���C��81W)�<Lt�s�ҿ�D�Gg^�>�0�9N�UJ�2~���ì(ôe�F�|԰�%s��Ǯb8p��6f�8�p���j�5چ�/��A�no�mi|l����w�?�ۯ������#1|$�����?R�Gz�H��#3|��%�Gv����G��Q����l��t��t�C�C'D&DgD>[�[�[?\>\�\�\?]>]�]�]�]�=�>y�>9�>y�>9�>y�EiQZ�-�y��y�	�C��9�#svxO��w��]�~���?>>�:���|�#6��뗭S)�"&s'�R�eL꾱6*�D2+�mJ�4��?6�5�O=<�ͶMm�w�����/����~i�����s�ٮkO �>?�����'j@*G��FdZ�!�K3s�X%��P�N�����2u!+���m����<�ri\��Z'i!��fd���͟��;�n��Y������g�S�ޔ���3�GR�{���L��Ɵ(��wؓ�{�{���Ao��4N�vq�O;r>:��N�E�KJֶS=�|���p\�� �}l�������k�~�s�y�q^ܓ0���է�O�N���v�~����)��~wO�V�_�o���I�>x}Z��X�O/?>������ջ&|���K����e]<�ǿm��z]oj�-�;Z,���&/��W��O�i�Jvw����n��ޚ;2ivO��TUah�Ed�ő�d��$��P�k�ֲ�L!D�Lc�;������o��Eg'���#�]�#�{K�=��(>�Þ�bNi҃�x":��w����O$o�%���N��d�GJ>��H$�}ħ=������g�;���фL��v���-�'���'����T�d8�G�S�{46�����ԩ�����~���^���Ȼ�Ļ8��-���k��eE�-$�dԨDg$
M��HTV�5D4�Y�����#2��H�I�;KF���tz�T�c��cߧ��	�5�J�ɏ7����ؐ5D����KR������{�H�v
喊������?�hO҂�%�M;�OC#X�Y���dRlY�EY��I*��$k8�I&�F4����u"�C��UD����b�U�_�KJ�������י&�ޙ	�T�*jC[�����r�#�uҘ&�U& �*2v�M�x�����ʞ>1�v�g� ����o�9��hD�أ��#��g�ݽle�t�2kS]�,�(�����%���2�Yܟ?���n�Vtvr��9;��?�!�iS'W�.u�m��4�����,��,���ɢQ�5���*�:Q��������H�3���n���Sr��5
�?�m���ڶ>����ܾ���?{��:�����C~���Lg{�:��\�紆�D�iե)#Y��*h���Ņ���$�l�[�|R���h�<�)�h�Ħ"�Dbߌ�͡�N�}��WǮUkxII~�aa�vFƚ&yK]/���Q���>v�$��oc���d��8US{gTBĐfh����2�kR|6�J��B��T��b�L�BYۤ�=��(�v[M������>9���	Y��~Y��=1��Wg��FG�P�������ك���~���O�����
����$-4�.��Ϗ��O\=���F�[�7������n
_Z���l�ߋ����ڟ�������\�kĔX�|�Tԛ��m��&�^&��=��C��#>B��,B�%qW?K����cH�F$U62&7$w�Ѥk���}�NX�`K�{�z��� ��S�I��W��Y�ᥙ�+X�f�΋ �j����ik��>�7.���6$�@[�o��}t*�<Nu[+����=:J(#N��{�jM\_J�����~�m��vk��ʛ��z��W�N���%%O~���k�$�0�61Fwm��RY��U���d��t��5��2uS�>b��$��p��br�͜��m[�;�V"m�-ֱ[`�3�19(�³;�F�1�K/M�'"eB�Z���Ϋ��>=o�7%2�����|���|���O��O�����&USY4��Ͽ;$�[�������q��%���˿��y~}�~���|�D߈�y�诛���������~�� �V�a�d�n����	ջ�q����i������^��h�g{��tB��_il��c��y��Xf������Kw[��M����ڊ�Пu!�\�KY��N+���D4yN�܌A�:�:���,�Y�p�'ʾ)=u���P�t 	޴���-R#ej�M&�C �f^���)q^)�5tGb�(������7y�G�Ǭk�2�xB�*@X�^�Z胴��i���c��H������:%ݚ��#�KL������d_�A���|�{}
n�)���/�"��4�� r�ǶQ�K�~i��d���6S���/	��-�$�*G��`l�K������t��ҷҩg�Z���$vo�SܻG���i�3m�%�$��B��>1ZX}G�9�O�9�T�ufK�u�E�N�H7yUM��J[��� ���%vQɸEH���T�t�������?|9���o6�yE���I7��(�ս̤�(�T�E#H���Ҹ̈́~J�&j��NEU&R���LHt4JRsȂ�z�;?�D{�>��;IB嚠���E�P-�A��ܻ�X��ɜ}�Ӥ���ѻ��Nv	w����zrY�]�^�')���&�{�_|A���o"!��|�b���>5"�]@;��BX�	�9)�I)�}�,�U�򺎈�M�<m��)��O��2$��b�d:�b�_Լ�'.컳��?�o���j���b{*������\��O�j�#���6�m���z�Ï���eL��nD��sg��2/��o��^������^�?�'��u&~�@������z�a�u�`>�����G��~�~�}�>:�޶�������ƭ�k���}P��H�������|�c��/>|X��F�6߹߷������{��������m���JȎ��֬����N�S��5���կ$|]A��8N렂$
�-H"� ���s��+"��C�����Lr��ĵ.sTD�"bB�HVD�y"�9���}��;0�������45�_!%$( :��da�C�'�ez���!����4*��4 �U`Χa9����6���p^&�CzI�!%��XBlX	��I����n3!����M�3��G�lPTC��X@4* �[*�+ ������k�v�0��]�h�] �c߄�H�)�UwGH�q�+c�hv[�X0i�ҁ�l�K�2i�����Za�Q{���mm�z�{aA��AN����o�f�vS5s��g;>�E��)?��B�wה�!�
���&(�ϋ�v/�[�f�PD���v����/��Ɯs���
T���TD�7����T@�n�sn���o�ǽV}V���V��&2����*w��Q.�;�P�s�9Ǹ��"�h����*.���L.�:Ğ��a��/{�F�4O �'��vD+�s�X@�ME�Hq�K����l�*݄�H��F��-��5��A;�1mw�Jq�D@�vS�=v�[ v��Wd����c:V�,��gSP����ڽ�
nֽu��c;V��Vl_@݅��o']�r�]���]��P�T[�6�N�M7�#�}��Op��4�}qC�}��V��f���Z�Cv��v��s�y�#*�k拊٪0!=р������R2�Y�h�y��f��`�z�)��d�Vr�&ⱀ�������y�y��v�����, ��T�{��ߡ�X0gs�Bl����1�;�M��܆z��l��3��,)�*y�J�Pwc)z���,i��Qn%X��[���$���H�za�G���@{o�-��Z"��E2�k�wA�T�0�vS���R�x*~�kF~����t�*}3�������Ӥ��4�w��w�����������{�Z>�]��Q�f]�NH��WP��fjauW��݈���5�G.au�� U6.lI�ʤ}y�G�K�ڂ��Ί��Qƞ�{�����f�Y���B!!n̂E
.�EH�cu����V��N�tV܋��52.eZfMH�������I%"�e�S�]�^Qsk��y{fCTD�&�YRD�i`	k�版�P��v��zV3��m�s����J�X\<�*Ic�3x�Iߞ�kg��e=Kl����
 Фa&Hh�X@�M��{U����Z�c��,�Z���%i^�A�v�����%���3�7���u7�Lx��Y�`�H�Ơ��a�<[h�C����. o��@d�{���ѷ��3P+_ƿ�[Ќn��qH��%uPR=4�U�- o�a]L�����_����E�ЌS� ����vh��<H%gm<�� ����m�Z�Ur�fyQ����,���¶hR�-���P,?�n)�=k�R�-����V��]�[��q5"�M (i��  g�ؗ8i�p=癗J�R"�[#U�D�·U�U �۝T)��.�<i�(:�-Lw@u,1&pҐ)N[�<z�.�XpfE�r 
�0�"�Ζ0ti CP�Ե�T�J���S�����\��X3϶Q˪B=OZ��F�3�/�OS�ԝ��:1�N���s�l<�p��t�3�f(���*���L`�˂p�ڂ��ϊgv��=���;e��x�C��`3�������ڐ�ߒ�04$�#4�,0��,�Y�X䃫9������"{������W{V3*bq���F)� +���P�&�������BW<�fp�659�f�2H����Zfy�/O����<�uQ�8lҰ|<�\�ZB[(�Y�.(�y�+oe�Y��(P�Y��N����K ?8m����?Ǣ�{��w��̓��ef�f�s6W��v�((�1�%�BC'�\Kly�/:Ů�����W����Oj�����rQ;�NW�u���m�|[o����ꝓ����������O��֟^�D}�u���PK   p��W�C��B	 )	 /   images/3fdb3be5-a051-4eb4-84dd-e907e6f5f8a3.png �@x��PNG

   IHDR   ~  "   ?f�   sRGB ���   gAMA  ���a   	pHYs  �  ��o�d  ��IDATx^��w�mI�؇��s]��Wϛ�~�O��n�����B�
 ��A�b($E0@R�)
@AA4��b�fvgvfwLۙ���~��{嫮9.3�G�u�^���
�A_��w�ܓ������?���.�c~Q��UH[ �B�sp8E	w�>�H������v�H�H��ʘ�n����.~|v��nD�lA��ʀV���.�*�?�2;��J��s��~��^�j���9�kg" �t !�����;̭��¸b��S.�z��_&8��23��ء:c�(ՠ,8��!��n2�dB��H�]��m��K���<Efڸ��s�!8$K'^aJ�dN]c��A��ߎ�A�u�Xa�� �@G	���zc�������rǈ� ��=�"���.��u��5V��k��k�ku_#׆���G:Ɨ>�����`L	8��H���t���ߤ�p].�g�GkR:���Z�I�h����i{�2�n=��Rcm��?e��+��7Oי�z�`eM�Yt����s���Y��M�s�#����ͫ���7��KoR%B���vx�<�6ϻ]��} 1y�Yi���U�����q�_��>��޿�<������V ܼz�}��ə7��`���Ť��X��]íeGs�>�~�K|���������
o��Oy����ƙWh%]ff�H�sp�V��L2{�i������?��m����9��/��?���g�����>w���;�u;�q�Gܴ �Z��Qj��!�j5-QÓ8�@H�[�x��H����/[�@E���a)��~�LYW���*.^����9~���.�_�	� �`�!A*�&��X�����X��嫜�x�s/r��5�\�Υ�W9{�.�����ܸN9XG�T�������=�_�ԉӼ���_�ڍ��� �H!w�j5��C���:P��{��5@���e���w��b8�:�T��~n��T�Б�f`*�E�)��K�!Q��V�%΂���`6+�C�SL.p��:q�����֎�B�=����_㹧�`���/p��Y7Í	��"ѕQ�]F�Ξi�#��#����L&a�n��GPz���&�:C�b�8��"�
�*�_�-���6ktkf��p�l@7o5�b���<H�,i�d��>��39������;��m���Glv=o�m�$��Q傪�c��!#G5�J �G�PP$���<K&#@	��������5��~tގ���J8Z��:A�
�n'٨;��TU���_�V!��+ng_[�>�����ۿ�'�z�K�W����Λ/�!_*��_��x��,��c�U1���;!y����V�.�/nR���"�J[ 8RH��ݗ!�Z�ɢ�Ack�d;�� \xQ��ݘ��^opb#f�\�O��O������9N����ߺ3�k�9�?�5����%��dFo��;q�����ދM�Fk��V�';�zE�F� �_Yu��\UV��q�\pf�l�q<y��yFH�4oJ����eV�[,6Y�*<�$+-�e�c���NЮ:UBV�Y�<φ[�������mft�.��k,'WY�\a�>K��9H*P֚���[c�\Ad5Z5�G�"i�ը�+�t�H)�����T�]�JG^��z67��y��[$ڙ�3KC*+�T]��湲�R;�? I�&1�#w'/�D�C���Q�V��DJ��!�$�4Rl-��\������}��X���0��pX�Ќ�)�{bһ:S	i�I1!�[�AjXk[�ۖ��c=�"ȵ�-%�I��:��iU��6�cr|�ɱq�'ۤwU4Y��-d�A�Д�c�a3�6Km�J۱�0TG4��Iǌ��3?��� c/�K!@:�(q#K�Z?Sc<0ϱ���� �B;)PZ�����EK� �� ���F�-� h��Zm�6
�^�4��L����E�V���~�!(��^@e�Q�f�"QJ�j6�#�8�4�t���G%�R
�5X&F:Ag*aϜb�XN�`��C�rĥ�	83�Μfq��7�J�Y�9�;Mc�T>����8�� ijf�79w�76�*N�9ޚ��iIR���<g�z4�?�L2�19��"I���B3aTPT�"��Da�ʊF��O?�����������?�	�fgPJiE��@+H(*E��0�(��l����$��ll���� Ǻz'o���Z���vgƘmǀ���2D�"V��Y+�A16:LUYF��EIQ�dE� ���"/ɋ���cQ`E�����"���f��4��ݱ�~����B8p�R&�?����1��4&ꆾ���a��E3٢?פ;	Y��A��U$��XE<�5�9|`�FQ����8)<�Y�k�:�`��(%y��C|�'��'��c�h4$eY��g�����
�t���Xg1��U���wο�c,�V$�B��xY��,�d�6&O����Ϩ*3<w�\'�"	��r��0�o�ɏ1���*i��X�&�4ҘF�E����� 8��+�|�g��(-9���ԁY�����Q�'��=3y���)[�����#L��9�#���.�퇌�
a%B�ʜbᰦ?-Y�'ω��
ϓ�
������I:���3\r�刴�Z� ˰�#��J��DZ39�bzj���ͦB���T�z}66�Xk�x�cM��H))��~?����%�A��nxL#JBC�Dҋ}������x�GM/:�W,�˅:�z��Dd�?��	��/���9z���/}������W���|���׾į��|�k_�k_�"_�ڗy��h���BQfḐP*â�b;���)f��LVir��ƴ)Q����Z���,)(&s��hf����݃�� �na5��Q&������2Iu��	AP�!�	�u����؞��K;���]@Q���f�A��ID��06Ѣ�n���R-�d�V'ejf���)ڭ&Q�Bx*6���~~jI�p#��-�
�UDak�lC�Σ@��#�JE
����.��Bi�7:���5��1�w�_������/��%��׾�7������o|����_�
��ēz�f���$��L���p�XT*i�E�����<#����:���9�qE���I����*M҈���3(
t����K�2H�0QN�Q��#��#	��#C)��X���>��?�~����}��{�"�\��?�_��G����O}�i��#�cy^P%�9��ȭKȭ����`��0
�Fk��jP�����!p��w[	L�7	q�UYˤ�8�4��8�V��(d����g����_�ؑ�9����q��>�����8zp/���s��u~�ƻ��np��>�ѧ8�w��z�7^y���f*cvo��tؕlWa3M���AHp��mjQ�A�@Z���:K�p�9H<S`.�(�Ѻk��C)�lQ�	�[ZUI1+�P�-*1����4�	+�������y⁧8xx��.�����~�C���������7����g�x�{���n!�d��$�?r����|���pב�\�v���n���	���^Q�_��X�?�pl)q�� 4Ҙ4���jx���$�?��
k����/�
k�.	`��(KLX�EYz�]kJ�zs�W~����]^~�M^}�]^y�m^�����w�����ƻ��2yVGqa��������������
�,��H�9��<"D�R��C&ण�s�A��6�
᰺�؂�.Ѩv�2i�W>)���$y��Z��F"1"'�KX1@#�A:2�E��N���s왝evf�v����3S읛f�����4�M�k�"M�&)�f�^%X�p���W����0'Ue��՘��w�R$i�V���V&!�.1�*�1^�P/�Z|(˭N}{��Z��\������'y���y�����8~�}�:q��~r����fqi	���y���;�F��_���ʉ5:{5�4�>��
Z��f�9��c�վ&v�������	�E����"���ӞUL�4�:���ķ�D�BG��`�dЏ�ES"'Ǒ�qVo��V
�Q<����V�7x��I�|�$�v���I��-�WWYXZFII�(�XX\�ҕ�\�v��K+\�q���<����2���e����C��8�R��!��*��o�2�RV^R�q7$��X*Sy&��(l8Z�hE%�A�l�DZE1�en�M�X[��¥���p��/���K��"�/\��K���Ξ����j����{y��8�� +�M~�Gʕ�<�t�ܾ6q�A�����fȊ! V�2����{ĸ%�ҭ.�V��W���7�t�K��Q-�0ln�2��#bmpV����QŚ�=�03A)��l,7(���ȃ�Ç����g9q�,k]nܸ��S����^����4���ӴZM��5��~�?�����Ox��wy��Y�׻(%BPUf��ڿ(Ҵ�)�]m��@��
p�M���y�T���?��	r���w�����XZ^aqy���eVo��t���n�Z����K�t�=����Ϋc�i堤�^Q�e��hҝ�`�5FOKzB��\[�1A���h��2�`��ו�8�F['�p'��Y��8���ĲA9ߡ?�җ�߮����i0�C͌#dJ�f�T=A�N��뼆NkE�?������7�����7���%���}��o��./����u^�]n-�`*�R^j����uA�R�F�(IwV�L����?̗I��j\�u"^48�`�1ȼ�=�� �q��X������M6���cL���&�	����#�9��]���>��s����a����zt�lV�ْ,�)ݎ �K��C���Y�7�%47���N�	w� �&���5��K}�[�Ča��)�uL8����FD6�X;8�ơ9��	j�X�Xr�JF��sH8&Ff�F��
)5�L��A9�~Q�s��c2*SQd�b��UR�ng7#�+��C�?�,�m���Aѓ�b{[v"��&ۍ4!I�e΅�h��A�_̷Չ#
��ze:��������8J���E`���T��.���ތh�ξ1�cஃ�c{���?�b��R���+ܼ�g#[&���K�H�<�i�:��q���.^Xg�z�VѢ35���0ձy�{0w��88A��`�$7��8sj��f����
��	��()���5eUqky��W�q��Un-m��HGh%��!�F��u�9���*���f���(�N*Q��J�!�9���7.0Z��_uC"!����,���ЁsP ���cK��bPR)8�V�\���ҹ��R�)-}�b3갩[t��"e�J��\����rN�o`�*ק�,UUQ����͛�z��F���\�����uM?�P6'(�q6U��*�����\�������U1��.H�ɫ���$�H���N���_z��|�eN��^�"�t�`����2:��*�^ex�@��2n��5��z'����	CY��$�xRU��ÅP�3[I/Jy:nZT�0��6II� ��m�z!;r�������[��_�s.l���=����ee�G���]�Y��g�ƀ����[�/lp��[ܼ�c0��8�"��-*�}��yE%J�|�lY�����z��k,-o�wK�AD�l�qq�՛9����pv���B:�2�L���>�������VVy��Y�y�4EQ�QJ����������ӷ9w�*�^��v�K>N`J�5��`�Vb��S`��b��wg_�;�2�3�sT�"04�W�����5�h���Q�$đW6���v`J��>h5
�����9K�4cz��ڋ�$-�hT��a��$7NL�v6�w>�{��湄�-V��Q�M�f��I��C)���&��h11�fb��D��Xw�t� �w=�#�aV[�]��{�,�s�D�͓3,�t�ؕI1I��`V�p�i��9��A�wTTdX��e���_��r��"W��d}}s�X�)@���~uM����Y)q�@)?�8@Yd\!�"\��jHhG�9���E
���Ғ�
�$���@';\%<�( RI�����*��M��~@Wի�vB ����}<���<8����go14j��)���2��G��T���ǙTS��Y����vt7���p`l���<��!��C�������s��;�޹9��t�C4Z��;6Á��v��G���]�.���a�ʈY�27q���L�{Ѓ9��������c2;;���:�O����ަ,��6��S)Ei�(B)�s�,��qL�Y��4�.KO�#�i4l��#�1D�8�s%;�鳁�u�
�E��DZ��8[�$�u�Bx2.�#%�
&���u�E�7���J:��8If��Z��;\���������$q̩3縵�N�,P�I�aSg-K�a�Y'1V�4HiЀq
c�Y��a��'V�0H,
���ʀ�% q6A�)+�� ��:�-i�0?3��Ch5�\�t����?����Kw3C/��ێ��J�'�7��̰��?ϭ���@!]к��S�2�%r��s�4��Z�e���V^`��n�8���	T�u�J8�tT֫��Rkq���%6 ^*���������ǟ�o����c����� Ú
��ZD!� �[s��r�pQY))��ʁu���;o`�B���B	�� �*H 
	Jc�GQX�8��%q��.^���w���?b����w"^H�	k��s'���
;�(<�%ֹ-�_8��Z��������V�m��	��V3EJI�?ڂwB��jg�^�TB����Y��vaU{�aG�UX8R%y���������ɉq���&t��o洄�"I���/8����X�H d�K�,�:��	��n�%��g��$�80���r�NDeq�{���H#y��W�����~�lv��ͯ1��I�`�"V�2�t*��y]@�٠�*����_e�*���	!h� ��`;�`Wī�"���k<��GZE�,/���*RJ��@b��R	қm�1��WIX�*�H4�_�"�����x��c��;M�a�RG%�� nj$`*KQ��ı�E3�#����Hy�}i)sC)t$�Q���đBE�~}���V�)enHZ�B�/�޿-H54�AU��74N8�o�q���^�LYn1�58'�ڡ��V`*��_�(�
�z����đ�X�A�Ee��o��ܒ(Fa;�=��nx1��ˡo� i����~FQVH�ͶZ)z�c�-5�o�%���r�s��YG�8�Hi0y�c�n0�z�7�R
��2��H���\憬W����@�U���'
� �T��юсjz%�:�혲0YE��#�$�Ғ~�@kIڌ2���cF��������.��aؠN�a��u^).����y����k�c�ܝ\Zw2w~0߫�=�y[��z}~�OEUjm�ɣ&P��a� �UB�#��&m�l'<��m�*���E�<�5��H�g'8P��4R{��/Yr�S+���~�-d��yw���eP�G�4Ғf�AY��p�qD#M��</��k� ���*Ɍ�<S�_ -] �+c�(��0T��Q�����qfq`��a.��3:����پ��Z��*�F�I���$ʟAvh^�)���K֏�c�И�ۢ�f�F��Wu2��W��Lι��c�k�����Ѓ����k�Z�Pv�[/��T�Cj��"����"0ᝅH)���WI�2#���8� �b����!�_\H �w�[t �5I����$đ�}th� �б��e�V��(��s�,*��W^J�$8}8K"K���R/�$
�!�����vֶOعR�P$��wh=i~��gx���^S-!<������ѿw�=��f�I���D�ƻ^�/�N&���ި��|�J��@%��|g�&w:�Ö2g�~��3.��6�o=��ci�Ń��(��"0,R��g��&h���V �B)�EEg��;:�HS�+X�L5bj+Y���E@)%ic�%/Kp�L�9������@z�EY��V����(� ��O����H~��\�S�eUy~�����HK��8HJ�y�DMe�<���g�P	�E"ꗉ�c��Xl��`�XS������o�dPRH/�S��4�]�s�:ܐzc)
������B��r��0��;G�Č������v�Om�#+*�WV���QV���`g,B�ЛPa|�G�uZ@�7v��8��`ye�n�OYV$I���F�ck��73��������5����mq��Zi��=34���'�j@I�͕��)mA�3�#��]'e�so�#()dK˫�z��KRQ�H)x�����sO����&���F1��KKVZ��Z���2?}�]n.1�i3�i���o#�B��F�8���G��y������:@��PV�W���_��wN�pk���I�8
Ɲ-ܹ��j5z�]�xw�/#��SJ/
���{g���>���3�� ����E�5{� Bl��֐۠VAzr'XY]�{/�HQ���=�s�0ӓ��H�}Ղ���A��a7;�H�������!�.\ac�KUU왝�C���/�3|��'94��$I��睠��ue���>��_�1���XZ^�=�d]ZQ�LL���C��׿�>��ط�{��%�C8GQU,�Z�����~��_|�յ�
�X�@�J��e
�c�_�Cp^�W��B|�"��ɭ6�^��=����>�̇��3�c,�d�Le�Ny2SkfF����+����Np��5��?�o)J��>�i�~�Q��#��5e�g[�B�]��X돍�����h�x����������������n�x�G���~�/~����3KQ�E鏚�
�Z�~��4%�"ʼ�7������ҏ����đ_��5i�̇?�W��)~��el�M��މ�l1��ZR@#M�:��K~����~�^y�k$I��q�`+A9��������1y�E��gv���v� t�}z�n�7������=��̴�{���V�\v��r�PDK�E/l��W�FID+i"%\�t����#�����~�g��s�3dwg����C�^���
�K	�fūc�u�9�8�^���7�y�����_��k�It�/}�3|�K��{�ɉqʲ�[�<�O�eiy�f�/�~&Hc����?��C|��s��~��8��y�ş�9���9y�<Ue���������~����g��Ǟ��h�����_��:���J+��E>������=���}���RV�O��w��{|�{�����h��[�7�m�J�԰^L�(��Nw����0d��$�8��g8���W��s��Ùdл�_5���uUɾ}�|���0;3>��St��9/����,����I��c�v��E ���K��j7���#<�нtZ-$ǁ�{y��{��?ç?�4��c��wy�G?�w��;�8u���i�PRQ�Bxn����X���?���nz�>���q�7��9{�2��9ȇ�z�������G���hpsy�?�����7�������CJI�֎,kh6.-r}a�O}��<p�1�x�*#Hӄ(\�~�+xL𤭑����3[V>�t1L�04���0��A*��_y�?���q��%�R�Z�-N�瀍�.�>�(���cr��0��Ƣ�feu����?�������.�V�+~�q�=�&mnv����gٷ�#�IR��쓏��_�4����L����z|�O��}��y�W����^]iԐ�# �r�MΝ�AYd8kx��x�����B��?���8w�"���3�گ|��?�!"�YYZ���������9/������G�~�k�̹K���E����3z���6�f�7��C�z���r�r�[���ʽm~t�o���5��Q���N���c��R�ҏ^�w����%�@��
�e��������{�������4�������������0�p�]wq����9���˜<}���5���e��N��f�lv{�>����y��G���`ei�wN��=�?�Q�'��p�o~�E~��k��E�4�ڭf���'��-�`�#`�\����:��f�봱β����F�_����'>L�$�>s�?�����?���=CUY����v����[Ͱ��dW�.�e�v�={��茡���ū��xe�/���gvֻĹ��Q�6~}�&���N�� 	������➱�;������'�?LF��~:'���ǯR^�q�~G4yQ�\��"� ����̲o��V�w���x����yk�$�贛4)�Ի�I)I��V3��HHS�����i��W��K�r��u�R��3��=3LN�qp��f�A6�7�᏾�^�]֖WoŴ�)i��H�Xi�h$4)i�$1�A�;���~��×���L�#��crr,d�؎0k|��0�g��m❟Tl�Z��� \s����o�'���A�$RZ>D�^qƂWly�o#MP!��m}�򉣈f#���8~X�J��*�~���/]当���z!I����vy<�
���'�?GG��m�ʫoq���1�gY����q��n�s��p��sT��nD�t����X��>y�q��3��,��^����ի<��k�����)sJ���Fa�w�c��%Rءo{�d�3������3I�Q���t��-�� �fJx/���IN���I���ҝ@J���X���Wy��	��6�2��"�s�9j��׶�(.�S����MмaX|V�AN�*�)�
�)?V}���CГx'VA��Ì;�V�_I�]���I����P��:RD���L�s��`�3x�3/r���E�v��!��$O�Q�*�@�~��k���Fc���}�H�N��E�$�����\h55�5qG��z�FnBIM�5q�H�!c�&�
aΣ�����&��V�E��g���S�{}��¨a2�z��T(����V�*(3A�Q��;>��;|����h���.eU1>�ހ�}���c��,ψTF�|����?�p����m�N`��ϋ���v�jY�|h}��Ј���~F�<|��СOm�M�;_w���H�$|РgC��<���&�S��	㝔v�I�ݢ�i09�0�i�n7�Ki7kfp;y�R��>�F�V+�E��d��29���4�4�KIc�ձ�"|d���R�0�X�08Y��>�TY��M��J�󉔵Wn���B�j8��y�dc��,�V�O�b���s����{��ػw��\��6�C�C5Qʇ��R���#��}x�����}9�����p����sϑY�O�j�(%�g�Ebѷ���N+E��29�a��I�><��C{8t`����=�}x�#�p��<��a�l�8N(MBYuU�' ���Hv#�$J�6��3����g��DIEA+2h饐4uh�����	"j�����^5RJ"�Ēj�C�� il�����m��lx���x����s��|�\��A�! ����sTe����f'x�����'>?�1����ʧ���x��=�$���S|����O}����}sM�Hb��7fYs��l��P�-����ŏ=�g>���ؓ|�c��O=�?�a>�����G�s���<p�]�M4�J�|on���A"�?�������cw��cO��sO�'���G�����ُ?ȳO=�ѻ�g|b!Y&(Kδal��,,�^IU�X35����g��g�#�=�'>|/~�>�ؽ|�#�����g�8q�]��/�D�8e� ��v*r�/x��M]�T1 �|/�VX�͚�F���1��Ǒ�{9�����9�����9��#�g8rp�sS��RW(>2�m���,R�N�s��<�����Y����)���ph�4��ajr�$�i�F��ɿj�FiIQ���������������G�ⱇ��ģw�����ܓ���c�s��w�n�#����������=����������C�=�O<�3O>��ϓ�˳O��sO�������$qR���w�}wg�?Y��8��^a ���EO]�o/
Eq�8� ���M._�ƙsgx��	��w���}�Sg�p��U�?{��'Np��./�b�_Q���Y�h�8'���nk-�n����p��Ϟ����$'O���s�={������{�q��M��F��q�������BI���rl��&�g���g~�^��晙�cϬ�>>6��������"�ٰ��H�� "����P�G���ga�=Ɓ�9f'g������Q����gn���Yf&����Q��*�`0�LA�"�0��A���$;�)�FL���"Ǐ����#���/��K/��K/��/���/��/��/������׮��}RmCvk7t	3��YƉ'y��y�����/��˯��K/��/����_��^╗^�칋�zR萈�*G�I"�@YX!eUPfL6 �sʢD%eQ��(�����Q��X+G���_Q/��Q> [a�>YY�U%��QEU���qk�Y誋��?�����]／b��3~ŹZ�����N�<�2��AV��8��	^x�5^x�G������k���������
���U^x���ɛܼrQh���p(a���e�Y���N�䕗_�}��
?y�U~��k�(\��~�O^}����5.^�H��Cɒ(��%[qi�UZ*�q��d��c�u6VX�u���֖o�_]dm�&+����Mn�\�9G�䅠
TR��B�A$�W9�����|����֖�.�-_#_��`e���E��o��r�l}	3X�U���@����y|̯�۵ �6�n;��p	!i�j�$IB�5A��=�W�TeUW��������`��9���d�v�M�4�v�;*�@�n7h�|v��\�EI����;����`@��b�7��m�/s�N�h�i$	�8��j�l(����
�"g�[a}�Uw��w�������66����Ho�K�7���N:-oe댵H)R
�F
B�HSZ��)*�(��m`���ؼ���u�7��������k�m�d=+ɍw`i7��(m���v=�����KL4�#0��-�ZhV;ڗ���(8{�2o�}������e�Ak�	����"�����$*Np*e��q���;}�w�;í�u�79{�*o?�{'ϰ����>���|��#H(�5s"fyu��'�����y��9��V�p��8�;'�����5y΁1�2�(����-{�ES�pe���aM%2��2v�7���8y��:��[��.\����s�4���6��Q��j��P�E����S�]�z��&E9�9/�t{N�>ǹ��x��)��1�v���><M:G�5��,[Og�:���d㩅 kk��p����������" �����j�pfh����2�[3(���`um��N���o����gY\Zgyu���/��;'x���l�^�_uq��aF��>8՜$nO��	e1�ʵ��y�4?y�g.����
g�^���^�ęs,.�l�"-9�g����VZ���|��n�l��J�f�Q��N�9�k�����Y^Yg}c�3g/������)�^����8�Ic��D�N��s��P�ѱ�R�em�Oo`�f��+�=�|�MN�:��Jw��?�2R]���G���ALy�E�F%��Te�}�TS�`��c�B��f�[�V�7�r�0X�E���)���+����l���Z�T3�IRS��� G
Ab�1��8�2���>yo�6ҵ��Av�����Li5#�Dc���,�-QByoWb������fć���|��1V�<�0(,7W3^}o��K�&Mb�eEY�A�������A?)I�`��y�=�?n� �HK�7r���ɥŜ�B�i��
6�9�~����!iU��`%�UC}�jL��JItb����JD��˳���.k�`����
�!�zM!v��S:E'-�u"$�~����k�v�A���*k�)�R�lE�]�*~�;��U:�N;�����XZ^�5b��������z�<��^	Z�������v�goŻ�� ++뎅�.�����7���ox�k�l��貼����&�X�5�y��N�[L��C���� +7�2V{�����.�=�wԬ�^�$��wY7�[����ʁ���U���NR�LZ�e�Z���!O
"��2��H�봘��n5�R��b��b|�C��@�Z�+��x�n�N� 7:L}�1iO*��	͆�;�n�w��aH��5`{�qE�!�P݁�?�mM�����.i(��#Ib�:m��:ð���q��f봈B�p��Ӥ�'2���u��pB��Mr!�dfz�����2�7N�P�3�4C�3��?����XEY:��'ݯo(���|F�zo�ؐ��'�X�_��v��P��m�,��;�ǯ��`i%e�+< ��!�} C�����3ت�*��u��V�7�8\��c�P�dC����|8y}n ��3��)}8��X[�se+Tp�-�2�����1Xg�1�;a���T�JG��#;_�c�3�Ae|�M)��Z���p$�p�GJ�d���ĉgJ66��ƍW cr�x��Jv���������7jTUE^8g�N�٘�r>���o�;�o�kIU
���Y
+�T8'������W�qX�ol2��^��n�Ax!�%��F����B�qF?R�$eFd*��^�n���v��4:ݽ��V�pX��-�L�:d\p�3p��'H�)|����(ۥ�
����w��8�*�kQ���h5Q3%m�D��*-�8��MڈH����J��2��8�VAW�m�?��8"iN5�<3I��&N�o���bI�*�8��s4ӈ�3m�L�2=1G�tH�6I��D-�-��R(Y���.ݬ���ĩB')I��H#$QlI[M�'s��ꭖ�С����H?�觕�Q؈�K=�6r�ܐ4q�}`hMη���3!��H�y����~&D�ֈw��u���np��!��O'��np��"뛛L���q�BJX�Qa*���8��U1+�m�Όq����t��:y�����cn~�,�^����~�1ݥ[t�x����D�ph)�Q�F���� �f����4͍҄>�//0=3���$���n,q�������&O?|���>ā=�>p��X���U�Ƣ�l���k7��+�YX�o~��G�15�ayq�ť5��>��M0=5F%#Ν����ר*K�
��6��3�#����|��0�I������q���r<��}LM��������Y�����
���D}'��Q�b7�� �+^�S�.L�}3S|�W>Ǉ�~�X*����}n-�� ˹��^�|�(s��)�����kPk�՛�x�g�^�љ�7��+��QV�W��3(*�z�Y�z�!z�]��?�=�W6�Z�̳�p���V���rV`4~��E������ￗ���_���Ν��?����ԇ�3}�^o�����_��-�W�Ɋ�Itg�hlWTHcH�/AV	�diL��S�"uvz�_��/��ӏq����9~�,���_繧cqe����?����B�ȤE��a����`K��#�LI�c���4$���_�G�ܥ+����M���/zg��'�>�{e�=��v��!GS�eQ��w��-ύ�ɔ�{���a�>v���&��8ki�[��?ϱ�G����9t������c�u�(w=Ʊcwq��]�;�x[ �%�1���sϱ�9��v�A��r`~����ÇHS��O���8侻����G��С����cǸ�c;v��=�ü8�f���s�=��8M��Ns��C9x���i��@����)�IA%|���U([���yv�)ؿw����Ё���uPJ�o~�{�>ʱÇ���"i�a!�4�59�+��I%p�R�c+��*�E�i�9�?G��ȁ}tB�����(
����}�Q�����(�`��c�XSEn}j�8򅉢Ȣu��DP��8!�0���S��{⚲�Vƻ*U>�DJA�|�^��N�Z")hFT�,�s��'�%TYEUT���T������V�/�P�H?����^�bR+��{�:�T
���]ai��o,�pk���\��̵[+ܸ��µ,\��ҲOb�Dڠu`�B���i���-"�9 ���(Y\^���nݼŭ[�,,����[K\]����7���������X�D��Q�y=�?��ʭ"7 �@~�^��/T<�_�M2��i�Y�Zl
]�mn�x��M~z�=^~�$/�s���y�w�>Ώ^?ë��˛o������3�vk@V�E�E"A���P4�b�|�L˕k79~�4?y�8/�}��>�O�x��o��{�ͫo��ǯ����oq��e�V���#~���A�������PqSW.\�W�᏾�S���o���>o����p�o�r��޾��f�U�����5^��EV�w**om��;�΋��G/��7��o�����7������O����^y��W�)^�g�	�r.|ա�zQ�r髀�D��j���7�2�
���k,�u9}�?y�4?y�4�['/�։�s�<��'.�ƻx��k�D�$"vm�H��gy��+�s�2��~���}��/���K�u�"o���;'�������E._]b�ϐ�D����1T��B�)�����Fƕ�U�^Z���.\�>��|��W9u��7WɊ�,���-�pDڋ�yVr��:�,r��"�/�
c,p��-._[���\�v���.EQW��c`8�m��T�[GHR(Z���]wg�23z��o����k��*׮/p��
g.�r��������M޻�ƕ[]����=�r��n狄�A�ss���K˼{�*�/\�ڍ�\����+������k��t�&'.�rkm�������:H#���_}%����@�K#[���_7��y�ZA��-{|�F���!�*�$"�}:�|�'kF��㘐�����wx�Hj��m��Č*p����D��Vev{��x�Dqy�pB��ȫ����f���jl����(�ע���Λ1�j�d�0�O������"�*So�|E~׎m�|굒D1�FL����E$�{4VQ���-������GA�Dó���2���ϓ�BU�4��B�����*��6wQ7
�u�k��!���>[�%Jm�Bh���O�-�T��\u֪(d������Xu6*c#*��o[{R���{Tܦ���.��el%�}䫱�j��{����Կ��d�u�6�twRɺ��*Q1�lލ4l�+��Y ��2x���&����FHw[Ф����P��C��;���(�q �l�'�m�> v&��:/�Y�;��Uݵ�p�g�;�|����!#�*�*F��V�la��m�T*AJO~�Vı����R�������.%�!����z��KC�v�nG��M���U���ͅZ:5��@6uc��;,P� K9�
�����o稜A�^u\�3{���2��ؒ�F!Q�DU������2w���@s7YZo�PE��~��y�q�������·;�0q�;��JKK,M�N��0o�thY�0��a�jg��ت,�����?:���A�V�$�٧�$�.$�We�O+��UԪr�Z`*�E�v��ϣS!uix�����!�ރ�E���/fUǡ<��W�[=����㹥�j ��o��6�4&�Z#��I�X�+ r��WQp���A�]�����'�P#A��������g�B?CyWaʑ���j�	J�l�y�<�8Ľ�� B9C�+�g��Śv��֡T����w�i�����;wp�<d�fPy͝O�r�vC������#���
�-��+*�MF�T�Gq�P�њ/�b�v���L���+'�ܝ-Zk���z{y�@�I�R)�.�LS�k��~��}I���F5�;�W���6:N@zFW��R�[뢈f�H�3F�@1җrm����!|zq��L}u���J�]B��+�zz�S��O��F�&]�B��<�C� �#2�@�;��-p��`BiA���I	[Ll�#�����P����w��ՠ@9�S�v:������t�^����@IK3*��VV	®ϲ�(��� �sT�2$p�7W������>6G��P%�ހ2D)�:yTg���yQ�n69t`/��w�6��m{b?M'>k���C���Y�r��g��Qg��2��>+�ޫt0�26�=VV����ү�m��l��=o�EbB@�r�T�O%2dd������u67{>e��f���u��~p;����z_������ֻ�\\aeu%<��C���2��ȣ��i���Y]������,oVr�5�� gum��n������sO���}��:
����+���orkq�,�i4�|�����|��Ǚ�gm}���M���?��[���?(������u�����|�����_�,���9���
k��yr�ד���:Zv�ɰ���	��v�,�Ɨ��)>��=r�Hk�;y����X����`fr�V����SSLM�16֦�j0=9���cc7�n��x���ǟanv��n�����pױ�8|� eex�ݓlt��8fvz���1Z���LM�351F'��OMM059��x�N���x�ٙ)�x�!�}�1��;\_�ŷ���/�=35ɞ��ϡ�%/2�W{�E����'y�PA�P�
�s�S|��O�W��i>��gIӔ+�x�����O����[LL��n���g~n��s�c��,�m/#�8
��"or���Qā�|����|�O|�i�֜=��S^{�8W��f '�}�B�~�gGp�M4�Z����YKYYN����G?D�tX\�$��4�LJa,�u�Z���n�T�?�%)ʒ���gf��IzU] ��QT%Sm������!�{}�&
%�r�M���'4�CR�T+��PYK#�y���i��Lѕ��w����p��u���<���$_��/s��!:���ƻﲸr+p�缓�s�F�9�o�=�8�������1���;?x���w���g/������,,,�7~�<��c����k_�"{�g�����ﱴ��Ӗfeni�%~!��Çx�'���|�G�)�Μ�;�{�����)T�h��ս�^��c#��x���n�G���������{�N���f�����?pe}��(h�j��Rb%1��l�왝FHť�E���?"�
>��O���bb�����yUm�0>9q\׻��KIԪZ)&��L��p��9�����������}�/}��|��'9�/eY��kos��Yn޼��6���.L���x��y��Rr��%�����֟��k?}�~?c�Ӣ�073�'>�$_����Ǟe~f��^�W�~����g�֒�Jo7�c��P2���<��}<���8�O����>?x�U�;}��(�����(ሄ�&x����
�#m�f���������y����Ad� B��U���#��9˥+����Q�����<���ؿ�{ʎP��㌎�����s�
�o?������>�q#Mx��G�k_����s9| �~V���AUVX����X��4�cm�M��w��e~����~����I��c%q� �)��Hk>�����E�����33�����a�ʧJ�4�ʱ����i�u�$������]Ν��ӓ�`�=��
�qvx�0�q��6�r�lqfK��%{���g��ؑc�����!����V�ԏ�[� �m�+�+��ױ�ࡻ��a�Ʀ�YW��s�;��|w΋�i�p�������ʵ���v������/}�/|��<�������YÛ�O�?{�����p}a�*�d��>���v:m��0_������>̓=p��=ʪ�������č�K�\(���ePT�2�+�k�P%��!�}��`�5W��K�s`�8��8J�F�B#��Ӗ��}ئn�,y������b�� M��Q����R*��.W��`��z/Y�6��<�����?�3O>�������Q��:L����]~��wx���y���()�ø����9G�? �#~�~>��'����l�	r(d��\�]�Iĭ�U~������[�z�I,����(�M����@=�G�(�E�n H!)��+9�[�ܱ�l��-pΗK�k��1����x�S߻wΡ�$�C�L�W�yC�j%��Ož�֝@�:0��ln�\@������D�ٹq��u��U�������U��.��0�H��H�"�cB��]�;j�����PV�i I|��</�c�N<���Y��{��IDQ�T�i�`��(ʡn?/J4%���+(��网>��U���p�F�c����$�)�4�W�n�D���|_����P�JBpP��R��;"1�s��� ����[�-�aH�^�BH_7��`t����"ԕ����k��!B�i��h�-=^��l6p��d�i�V~Ui�H�����X7�N��h5>R&ˇ9wz��D���+#*��s���(}B�VӧF�c��-�DZ��:�	c�c�R�e>h������޿,�����E3�/�����9�����JU�?+{r��c߬�;S ���ɫ�{r�Qjm�=��̴!a�j�|�ݎ6?cL�:)}��޿|�7��d��k�,�}li�Fw�����Dn��}�k?����m�5s��F
�k�EA���Q�M�Uv��@��z����7�Zm����0:�^�,��9�7�'�gƘ�q�7�e���G&DA�}U�*(|j�ŗ'�!xs/��"|f�`���>�Y_d�:o���T��2]�QJ�Ԗִ�.�'τ�wkS��֘�=�c��G�DK���Lx�e��u�ۥ��_�QD(�XV[q����Z�H��
5[�ڹ��I�dh
�'MH�b0�6�!��ngy^R��f#�2�<�}��Y��mj$�/�8��i�s^�;���8"�#��4�0���H�m���Z{��J�ބ�M�a�DҒ���Ҕ�ǃ�ć�V�*xtj�����	1��'��q�뎣�˕U�m�5?PV�Y&��V��a�}�1e�$s������s���R�P�P
_%˺�Ӷ�����>��n�y??I^����W�k|e,�%N�lS;�n-���|����񒬬@i�ʫ��4f-%:��o���?���Ī�7�"x��1�����B��f@��#Fj��@Lk��N#M(KɳE�����>fT�_#^��{_��g��>�޹Y�HS�>���w�����9���2���?ݡͿ�u��X��X���1]�g���;�{�����ݹ������m�|�
�G4�6?��}�v��6�9�t��p����o���7����i����)�$%����������v��z�X��K��Is�c`T���A�ȭ�J�9��GՈ� Q>!�T]!~sv[F�]/���
��j��W��kؿ���.D��+K޶���h�������5���!�$IS�9�޹Y\e�����_��h�I (1\���[g}��[�f����mh�%,�*�z����Gweh��B�P���o�쟰Hº��c���|�L�f���ͯ�[��e�:�;�����]�/uɊ�dA���s��c���}�O<�4�~�������;*M
I�UiR(�՜�̒s���q���ViL/���6~#:��BII����d�>e���1R������n��]Eܴ�JP|ć:u�FR�k��z��������_�*{���'��s����p��� �A�Z�m���;Y��5�q����_����Wi�)����?�?��-���&b��Z�t���L��i�>�K/+���H�7@�-D�uif�;L�w��&��+�ZZ�,j��W���znf�ٙ	���Y�����O��N&���D31�dnf�4�X^Yay��z7��Q��o�[�������O�{��?�D~��y��lX5U�7jJi�=��]����W��o�*�V����?�?�/FH��3u��L��<���g=�����Wx��,.-o����bj�ç������0�>u�wN�du�GY������7O>zG������'�^���Y^Y�ʈ ee�3;ƣ��{�1�jp��%�<q�w���:���l6�������o|���������?�m^_c�q��كH��f��gKWI7/pt�����7���č����?�?�/�����N-�1T���c���ٿg���1�:���)��fn�3���$��c�[Ҹ�s֍첰Ai5{f��۷�ٙ)ZM�L����!eDژ`~n����ә:�NǽV/�(���d�������La1y�f��~����f���l3��s����h��>�m�?�1x}@�WJ�!��=�A�!E	K$�pF��"6x�h*$v芽 �Ar��������J���K;A�X�,���q�`�
[X�am�-Jli�oE�59��e�-��6e����W�)*��=u_e��p�gQ�e��6��P��)F�Twh��3��[Nq^~��m�]~%������V�����#��\7�ZYgm}�l�y�ݠ>g�{k,n���el�E߻0m���Ĭ�������"�+�l &��p*p���7X^Yb������|c�{=���Ŏ����4iP��G43G�PxQ�r��"�F�1Ri���#R��_�:���Hsd���Q
���@�X�~�$F�m����Ϣ5�nU~��DH��*� @��� �ȷA
���4B�Z�B	�P[[}���4��+��ֹ~�2׮]gy}���:�G!�IC���Ƶ+׸vc!$�����6Ȳ����\����Kld��zDnǻ g0y��7or��U�5��n�[
o��&��$�	\C��h���>�T�,#A����S�wW.b\�ٻh���{�qy��o���(\�*���{e #m�v��R8a ��t�ߠ��3�r�{�e�5�����Q��;���_T��r���,�,�1��:�(��*RD�"d�-����L�e!�g� �?YYU�z=�W�Y���/fG�a砪���`emm�:����%���5s�.�qE(+*2����	e�4�*V�8��5�H@��,���4��8Ql���kB��H1���.KqY\��SL��T��}���3R\�=�Ȱ�&y�q>:���٭[�!~7ɦ�	h���I���!9�Fa��yE�+i�:L�N���Q�`8?p��:��bb�I#�g���@*D�265���&J(wD��sPY�ٍ�9�":}D�#��S\�V �@6�����B����J-}�\���Sp+t�+P��*	mb��c\���yĩD��{� �u�(�����*�uh]������z�9�O��X�-�{V������/z�d�5H%I�M�g瘝�a��B+�����T���j3;3���4�4��v�p�1��������$�T���1�~�
��LLL2�gis��z�v���F;xW| ��6�\�)q��ғ��+kq�3W�T����14
�T���an;?�ݖ��	�y�pE���A���{<��H�E }�������x��$x�5��t:"j����c����-��v;x�y�h0=1Ɂ�Yƚ͡re���|�bM��anz����F)�6�����gz�N{�8�A�;�E�L���~�y��k��P���*+i��}�eYar������AnY���c���p��U]�aG��f�0��V9�9�HLVa]�h��d�����D���*�d�"�sho�Yaa�;�z��<�m�d
��4�Mtܡc>��9l�ë?^��J'	��$I[$:%�������)�fL��j�RJ��b����"�e9e��1���F�}��Z�P#A�o�Wm���@��c��p8����nXp�#i[H�ïD�!�=�4��w�J"�@��J��L(2�D��?�	�l�7�C�@��]6He�Db��HT py��J �$F�З���!�Ȑ���Rb�-�!�܎3�U�`У7��2�_]+G�V%��O<`�ʂ� c�ߧ4%��W�E)E���nN�ʒ^�G�?��*�-���#%���0�x�EIУ�{`���;w���ѫN���WB��L����FT!���y�B̺� "��a5T��;/BU1��}:�(E���6�\���G�t�A�(b�w��R�B�ID���r�Ă��A�u7��§>�v2w��tZZ��@����u�^8ϵ�g��.�M�R�䘤�T4tI���lh"����¥�W9w�<��(m�x�1َi6L4S-I��`�[�^_�¥�\_�N�ۣ�-�M��`�1ݒ�M��h�l�����s�;��[W��&�-A���W/\�PC7a��F�85 '��QZ2F�;�,A�)vP�%�(�	l?�n�ԥ$M��BT�*0�
[ZP��!^\3y�1��E$%�l���^��)�KW1���C�3.�����Sy�"�� �U�����H}X���s�������dmy�3��p��9֖�iD�����T2ъ�lGL6a�)hh���"g�^���sl��"���鱈��c�)o*���Mn]�ӧ�t�"��MZ�df"a�cMkJ��4]��-q��9N�>��͛�2����uۨz�"n3�8�8�ɱ3`e�m�q���Wh\�U�RId��̋b��y�*��ܴ� �.�kYQ���1N�تAUŔVa��? e���q�M8+}߀��#�ҸR���Z��=T��
.,��v�u�-p��T'	8Co}��/q���7z4���vJSK:�������a"u4�d}e����r��u��Y1ފ�hk&ҊF"h4$�.7ظ�����q�:e�G)&;	���8�D1�04eN��r��u.]������H����Q,�;�� ���F�c�:����<���a%�߂<���42����	KNNY�SK��x#G��B�)Q���I����*��Ґr�B`(E�EG��D�.K�����������|���R��p+C@z��2<�Í:�-��6r�*plB��Bi�����G�IR�6�q�#'%N��1*H=�ykgS)���FG
�AE �"�~���k!���vWD��&�P>A!#LQb�M/RI��r���lt���f��<������_}����iٷ��q�gƮ1�h�l�[I�Yl�#����T[z	[��;Ő��x�U��N��Ѻ	o��@�e��wr���_C���}��O��_���p����Ks�P�b�}5���J�p�H�#���/R*��G�y>Z�3*]z� I陱"F!��D����Y�˽jW!��y���)uE�ʜ����xz_��Uf�st�O0�y�9w��;k<3_��|�CS}5�ĺONH_j��tq`�D�S>�YI��ڗ��w��}��C���"�~�l����j��E'��>+�ǡ�[9Y��x��.F�!8�����^ᐱ�$UV�� ��m�d7�u[�A꙯F���:��s��r�
_>x����(�u��G�p��ksߡi�x�&_;r���-�grӬ<^�([ᙨ��H�ʛ$�I���R��R����ٰ͇�>��ρ �C�k� �����(BAi��o�V��x��D�,���E}D�#�
U6pY�Hso�\e���Kh�M���|f���ބ��V�3�"%�ms��}������	̓�1_���U��=L��|�%��p� ����)�ED�[���ֻF�I�n
��s��z�L��߿@ �� �)(��0^/P3r$�6a��/���8r���2�r���j[�JFU�Ҋ#���L���̎7��}���8B�p&+ye镆�Hd�23��I��̀��t�%X����+㥌��U����FYDT b/&�
" �>_oC�.�-q�M�/8��.`�����F4c@?��L��/��n��*aX�ț9�o��=g�{l@E��0u�@S���
�
Jk����!�K��Q�-��[|�S�h���8'!.�c]�T�n �2�qr�Vb7Z�|��k#���H�"�s��Ų-����2yw�gJw�v�g<q6��#E�q�4�T��3f� �qw���>wMZ��׋��#	=�^�w�A�)�&��P��B�UđT��D�34���
>ɪ��C����k.�z�;m�@�v��*��$80�.���_DR?
B����!��i��?V���q)d��DT!ZB��K �R��=iI��)J���c�};��+6�Yd�@a-��������b�QP�����x�����m6.A��`�� >�H�I�6B*���{t�"�3W9RY��>��w�	���A�m?�̔��.*� lY���!� eR"�
�Njƚ��	_��w8��!P�$����bBj����_���A��)�%M��$�0���a���![����|����T�����4�/!��m�/*�ᑽ��k��H3Nx��hD\�wj$.�Y�H���Ѥ���X�Nb
kqB��.��]I!��&�$%8��ĵ�!��^���!�$�`s�\�%��#����\ɖ=߉�{���a�n����w�P���N�� �CF���|*s��!���HsQ�q�	�T��TY��+<��c��Y������O9LU������hR���R���*�BO����$���E�/k����������N��r��U�Zg�p�3�z��{���|��J�u|G{|���_�J��$X���s2O�Dӭ�\_���t�s�s��%Ξ;��s��p��.\��s�9{��oP�}��R�l�D�]�����9w��/^����;��.s��Ο?Ʌ��,=�c�S�+��\j�C x�R8�v1��0D��>��Np�w���ϑ�w�NR�=~�.��<�Հ��[y[��ad*�,�1'KN�z��'Np����>�'O�뿟>É�xｓ\�r�2��u������>�>'N���Ӽ�'O����S�~�,�O����w9��ȍA�]����M��-vʧ��:�h����G�m o��Cq.J}��p�A8���W�����P�v1�(qR_3w����p[��C�(3d���N�}���ϱp��7Y\����:7�_��,޸ŭkt�7��r�H�=n-���.�`�����׮r��2˷z�+K��M�쩃���"�c]�Ͷ\�Yxο �w.�2�4
�u�A⌥!��4#`�=~�K.�G�x�+>����Z�-X�R�$!���<����P�_SZ{zp/���@9�F+�V*�|�4��7�)�ek;�Y<S��}��B8�����nW�װ������h���F�Q�֋s����4����g�W�(T�^��0�w�rE��l�U8[a���5� �����c�ٳ/{�γw�>�<Ⱦ���?�����1>58l��!5�M��w�~���Ǿ�8p���an~7y/�h�7�e����6[�*��Se���9H�.g�?���}��H����	�t-ȭ&ڲ=WGN8�Ln�Gk��u��"�=�=��E8*]g|6�{�������呇�������������y�Z�J,�V�Áx��y��y�A���{�����㑇���{�����ٗ�GL3D���
l�=���8Ub�uP�w�t���j��م��������#��E���_6����i�'�� 8�+p��Ε���#	��#B� �"n5���a��<���e��}�߷�}{�ٿo�����}LOO%1/w'i���4���e��}�߿7�	��������39�n$�a��&�� .�s�uX[`�g@ET��p�jZ��};��|���e�2�u��A�-���B|���_/8Ƌ�C�S��߸��9փ�`�[�B!�"�M�-�s��2/ Gi�fP>L�L��HZr!�z9���\�k�s��Ob��!hR���ZPs��7ǼRj�`7��]��g�t��Ͷ��U���UVb몊мSs��W�"��2��2�?+�`0`sc�����>Un�*�KD�~��@����n��H�z�G��3hyP�O63^�����<�b��@�Tu�� �ESˣ{ӓ�-f��-D�Rk����A�Ǫ��-�Q;REH�]����"QZ��r�h����L���8#p���ܰeQ���X[[c}c�nw���{ן]'�_�z�l�lkr���x7H���w��
�QEYW��RV�ـw�W��쎽��9�"r���/;�pH`�,��Xݴ\\u�f9��ە�"�p�)��DJ���"�D.�^��3������[�n��ۏ���ZK�e>+tYRUy��l��[��� ��cKGC�4F�4�gM:D�Iߓ���x����hn>8����������5��� ����K�S��M�4p§W��g�p��b����q^�<�z���D�޶��u֯Vm`�M��Z2S*��q��R�:�5��������9*�s�{{�?ۊ�3���֟����tu�."�����}J ,�
�k�F��eI��,�H�74��}�ɭ>XWIH� �f��.<�P�$ZKb)�86�72N,*�gM�Ȣ�{�*�R�x��p�L�}�.��N0��w��x/ΉmnL�VJ
O"ep�vl�c����?|/�e6b0b�!iv'�;�&�� �vn�@�
!|��h�!*���r������$YD@SB�RR��r�*��&ъD8z�����s.�ȈM�n�!t��BE12��o��M����Θ�#��Ysg�;M{�>ON�6HӔ8���i���t���(��*�ȱ��#'U�!��VAK�u|�'��f�H��.�F�����޿�9F{T>�@`�c�����/^npu��Z�OVY�TĲ"�De]P�G$bi�LF�����&/^O�����,E�FG��E�\ �o�p)�4*T�rY����NI�v���wS�4	�d]�W�$	�F�f�I�բ�n�j��t�'$����z��//���;�����UB�P��b���VՂ���;B�w| �E��]��D%!Y�-*�т�XjO�A��*ί5xc����Β��u�Z/��z.��lQ��~�X�R.mXN.W�}^[Hyw}���D$�p"��H³�[�"_�\��|���}v��+b;s��jT�!��'1cc&&�i��h-}Ƭ`�l��b*C���>U�Gz�P��5�27��"p���P���Q�23T�g�Td�u��49
"�,o��9�ú&7�$�fO��:cF0��:(2�W��2��������|�r�w�/pa�q�=ʭ�٘=@�t8�:��{��k-���1~����^Db2$^Ic�Z�>�GK�$n����NcT)��H��o��*Kt�213��Ç�w� ��i���2C��lf��n�҆a5�B'L����CL�B�mzE�f?cs`���}�f?�_��������MM������ߛ96{��t��}8x� �338��2_Qb��kJr'*"R�\�=�@��$/
!c�I���?cT#�$�e�b/�ʺ�ͥqN������~����\��Lo��nZ..�,l6Y.
#�_cȨ�z�
�����F�DI�7�w|�pe0M�
b��a�x�Q��֠(Q�s����r��{hML�90�Z�Y�)V7+��\[.X�I[8v�~�#��Gܞd�_�����iX�+�7JV736+�����w/<|{ �MVz%K�9+=�Jױ����֣���w�{/�|�A��E��2�bK�a-o��0�2�Hb�Е1BZ����is��*�N���� ���4)PiN��c+ǩ�{�eYv�w��s�}6�͈H�MU��@�"� A��H�)�2=�Zӭ鵤����FK�%�Z�tS҈N� A� S�ʠ|Uz��6|�sן3ι/"��
 �=�f�z�/�{�c��g����d����;H����Fx?W���6�]�j�H�S�!~����.4E����(�>�SC��� {&��i���sm<��Z�@�iI7�P�J�>���S�ۨT�Iu�N�)םB7s�F��kA�ѡqf&��>9@5�e>�<��h���n*��I��5Ɔ���`th��_��8,�2:�Ȭ��O;P8��;Ǉ�55�@s����.�e�f��ߤI��Eb�!�%�!�UC���{*�v���ћI�ʀ5Ui\�}�xH�Cka�&��h��d.�{����BG�I�,�?��Ł�0<�������'��	*9f{�^� U�>.w�!W
����T� P8dʐ�g��Raҙ ���5�u)
�L9��yfH9䅃tB°N%���)B�b�J��9y�ɵC����*���z�F�sB�)�җ�kԿ�h�����B~w��ٟ
)��̇\��˂a�Ar���N��q���C����t��A��f�`���I��
-�4��'��#i2��Z�Y#�q�$iJ�P��a�ocLP����ݴKG�IJ����r�U��
�`�}�4#�����+��A��\3R��d�VV��St�F��,W[Dؾ��I����gN��DĈf!@��9�Ъ�HOUߪB^�d��r��
ȣEd@�n�nP�SmI��'/�0�Mԏ��@�w[ʑ�=�>� ��F^�-E[��3i��~I��e�#�,q��u���H�Y5�΋~�J�R�V����2KK+dI�����WR��i������ҋ#%Z���g{�HcVח���@;�Ȋ�x{~���4i��Q��n
��Oj�i�X��Q׹IN���S�XQ��&QQ��8�2G�mpMf��i��{aA�hT� ����
?�H��<2����g���NO��8�`*��vVu�!ꃂ4w�b�X_%wV�u��k뤅�!��7f�3�m�[,//���J�D�N���)~ I�6ˋ7YY]�ۋL&�=�
�F������Z��\�!ŝ*�n�����/�ٟ?C�
�=����cP�98*/L�#�-�M�NB��{D�#<a`��x�P8
E�&-M�u���� �H\D\ar��#{C~�
�<4������C5�0Ѩ�UT��X��'G�0��w.Kz����Ε��8�M��^u-׻I��:�̤��Q���!KS�L��u���VE�&OzdiFk�C�۳�ޣ����	�6Y��'�Z�Ϡe�gU��%M�"4:uQ�D(�uJ�3���T �c_@a���F��p�%�IA��"ÍN��8!�]7�Ūc�$��HZ~Z��Q������;<6���T�H5�ȶ�3PsȲ�<�*Gjd���z��fz���z������{̭Tb�1���@8H��W/ZY�6p}j�&́����S����Je,�0�ި�hR�X����Z��Ѭ�m�u���J���^�H�NCoF�s�̵B{�a�T
�H��rs�,(�F�]�9�h���Q��b�F��~���q���RaX,1�l�{.��#l�)I�s��6;�n�ʐ';6�7������
�ζ��x'P��f�ľ�?�������f��܆_A8'Ó��$)��T�*��Ln�at|�J%,��[On(P�*�� cc��ncxd�|zOH�FK�*LON�{n����?^a���G��x<Ƹ���݅6��4Gh���F��J'��d��b��G\d�"3X=W��UCf`��H���7��D��0Yd���Ln�5��`)�H��Q.I��C+Y"/RQ�ň �����J�s�2���\KS�ю�R��ȌZ ��!j�����E�$��#S�'|<�C
I=�V���=��U���t7Õ�CÌ5�4-_���[���6G���l����q�I��v�ב�D���S
ǖ=��&�ٺRQծ"�*NŐ��>�"��	����G��M+&��Pn�heþ�.n5%/��͔�/lp��m�n�D����+�ڹ
����K�dG��~��w�z���*�׏��"'�R�"'�3��Pn)�2�i��JG���,7��43��{ݔV_~n��,d�нGCX�U�ENRdh�"؂��Z?W�?�4��
rca�;���Q$|�>-	"G�ĸs56g}��(4B*r
2���Ɵ!���Jl\��L�C�OM" �FJC�zc-�+m�yb��tx�|���l���]b
W�anʉ�ᮀ���9�V��V�\=͍��n�s��2�-E�[����7���]n�-s��WZ���E����67ns��7V�I�h���K�,fc�67o^�ƭk�:�d��+�`[�ĝ�4��=��6��ϐ�.J%�q�b�٧Pfn��nߐҪ���$���Іw�eT�� �1����� w͞�O!w�26��B'�_���7��{��?\�w��ʹ�m�kH�E52�{��VQ*�P,Z�S��%g������lIB
�n���
W�/qka�n/BY��<l�4�yA�qsa����,.���E��E�
���,cy�ŕ+\����z�$�(����ᛦ�=��\�ڍe�W�ĉ��	�=��;ı#�hT�t�
��q� �@n�9CZ�!C$!B�H�A��qQ�Z��C����E �H]ҟ9H�3��k���,���u��u�`��B��'��!<aL.Q����&)@;׷�+���7��@
��~��t%�#{9�o/��q�����;�4eHS8����Z-.]��+o\��SWXX\"M3C�)7;]A���v9}���s���/���L�u?�8�4���^}�2o�s��W����a��a�Tqk��ۧ���9s�6�k];�77�R���&W�B)\!�g
�� h��W��N5*�Q��Ό�G�&7�-�K�#�9�7^��!rkH�uL��+�g[�)��dnJ���������~�p]�ѱ�N�����i�Qd���V���a��LC;՞��+3�r�&{VY��5�	D
�0b�r��P�r֑��&�}��#�S[���SH�U���6�_��y~�0�y�Z��_����s?�YF''�ï~������tc��;F:q�!!ڿ��-��V�|������V�!��aM��k�\��)[~�����SA�p����g��?�Y~��?E�^�7��5~��k���G����\����`K)�5�"�s0HO��"5X���	V�BQhA����=|�#IR�����"�����(N����6�K��Y�V�K?�S��O�S3�x�W����?s��e�: 9�v���v�tI-\k l����IЙQ��3c����
L���Ƙ66�"��5]�^�ߔ״7t�1E�(���xO�%W_u�t��s?�Q>������_����W�ȮǵcaFw4l)����BHM�uL�=�z�h�,��)q������Rj�Z5���Y~����;�v��{�V���%�9
����8U(lQ�*1/�n��5�.�m�>�]��:Õ����n:���
��˕B�
B�P��kjip􎊌*�S8���bмy����$EH���A>v��{w������?���1��qm�l�	d�+q�R(�F���%p2�ĹA��� p|��i�DB�(�3�t 4^hΙ��̚�U4Z�:x���}-yj@�[ˈ+<�W+����S����8�� ,��gE�J!5� C@ >� �c�O]ؙ(�{k�he����Jۍci0i��3+�%R� �;ᙙ��ﭳE��vߣY�Vs�{�Ih�֒B�8xA���&a`�����!��˭oUPqr\Y��<r-�����V�}������FS�C����������"%Cړ��5N%%���᰹ܘ�
��p�� DS�Wfܙ��Z	��?�Y��O3><B%��`�;H
�>Z`:DYץ��4� Mck�+���{��g��\غ=�*Xؑ�({���oy_�,j�^Sc�	���㞔ś[�2�lRI����w~�k������x�v)��?��Y�+���8���B�1���>�(AkM%�{����|��kV)E�$���o+A���AV�$iB�8r����� ���g?�8O=� M?ĕwg����?��0����-�u/�{�W��5-g��L��$Iy��|���{�����u��[��<7{��(p]����4Y�#��u��-���gQUܷ�M9��uw�+��-�����Q�,�q]�5�T�(]P$�P�{9��LL����x�i�����^g�R�6Œ�,%K⻬�?�h�t�����9��P9i�����Z�ɂ���=
����^XB��~B���1��g�Ygr|�J%xoE�?���[Y]ciy�N�GQ��Y(��84���� ��9?H��8�C�"Mc�~��F�S�XouȲl����}���w�6Ǒ]���K�O�[f��f�q��6�'�4Ε<�lN�k�)Zk�<�P'�V*T+�3{�u���g?�g�>;C�%����8�iɖj67/��DXp)�k|��x�;��7����J08Pgm���8�ݽ��|�Y>��#v��y�2���Q'](KX �4'I3*�������a~�6*�ނ8I�Z�(!�=<ϥ׋�RR	}�$%�r� Uh|�evz�=���k�\ǥ��@1�e5�t=�����<q�7IzƩU���@���I������ ?��#B�*�u{���YN��H�AJ�h׭V�R��(�17ʳO>���K�����Q*3�8mp��v�v��J��Ƭ���z4��;_�?�����[�Z21:ĭ�e��������<���O!�F��Z�B�C�H���B�c����Ek��|��������s��%�DѨ�PZ�$)a�#� �|߀@��t|h;>ˌo!I2�������ӏ񡧞!� ��ր���w����t���,����[�����]Z�=�[�,˙���ч���8�wn'�d�t�;D�Y��4IY[]�_�_��t�=�2����̅{Q̞ݳ|�#O�����3�c��HXYZ���1 �-s-��@�`��-� �Q8��v��מ��N������A�WB�o�v>�?ʧ?�a�,PEAQh��F��s8&�����`���&���������⍷O�nw�V+��C.!X��n�B��~�I~��>��>�1\� |�K�����?�|��/���N�{!��z�߳�O�i��/�,s��w��O$i��p{�_�Ͽͯ���pk]@��Eջ�&�36Vv�M�<�����ssS\���Ͽ�;'ϙ��r���W�;ދ2�d)���뷹|�:��PZS	�(F�����b��Y<7A)Hs��B���.0�v=Ix�Z=�`dh��{�g�~�F�ƫ�������7�9K܋n��p6��岯�v�VW�jw�}��|�	��O���|�r�\���˷�E	���7a��v�ϑ,,.��U�>y�N�g
1
H����a�?�����m�&N�{��Q�p�]��f���R�U�6����ͯ�y}U@�VA��z\KG�W��i���N��=����_�65�˯�ο���:�x�%�2���9�]n�Қ8u�}�uH����	�c4F�)���&(m�y�c��q����!�z�,m��9�#������?����������8u��4�����[�-[�~�������{O=�0�'?͟��aay���:��/���A`#�\���-�\���h����\�z���V?}����24�dnj�F�qGJX���e�M,��TC����O��{vq��<��7�_��YZ�@��q�ó�$���A�G:T�>;�3O<N�^��y��қ�=w�l�t�P��2���D��݉,�>�ex�VC<�#�7[�P�2�}��(Qt�f��H�f�ҦTy���������GiԹq{��=�<���t)pȕ�n�U��kT&6��5�ṯM=.H��q���Ʊ��8rp�n-���o�?�&�8�����|�׮�������s��<���z�:.]������\�v����E���f�,j%�u��X���y�^������v���^g��M�o����y��0׼z���r��5�ݺI/����cl��F�������o�L9W����TQRn�dF��&pS��"Zl��x9�f�Ya��f�M38P'1:m����m�N����6�n�n'"��:��ctt�ٙ�ǛT��1p�<7�yn�����n�@���(;蔍�h�|P�@��G��@�[�ĵ~](�4�����thw:�;�Y�7Zl����-�7ڴ;������I����]S��%2]'Z�No�:�����tW���8����o^`��Y���5ɑ��8�g����<OX�h��Ѣ�6�i�;t:=�݄<��aK�y�����)�ݝm	��ع�{}̺�۶za3�����#����욛��F��2��*+�/�D�Ȼ���k�Zk$�%�nx��=������9�Gx����=���nE����^�.0�@�}�<��A�
�N�0!e�l
ar	�k��88�1R}GR}��F�f��@�N�V��=j�
�z� �!�:�=;F��'�g�Y~���s�����Y�D{�"ݥ�t�.�Y�D�v7]��V��"c��L�y��~�1�S��T����V*4�Z��Zϱ������%�s�̂=���O�$�}��LR��'�9+>H�6^�Qe��q��ţ�����i*�O����:^ �-��� �B����;˴6ZTܜ���<��<td?#|��/E P��^��'uaҰ��R|kӻ�$�T݌б�o�֧=i��Z�E9Yd>B��&�P���N1�a��RH)��j�u*�*R�������M�e��d�T�H3�*M��o�}�{+�d	���w3|��C��)[\�V����+f��8!�J�����FkH)Qy�.�����#�$!�b(z���.R�$����z���#��4����>���&�Zi�<�P����:�lU��:u`:��MV����h��
T_u�J;�iE �,p�5��x�XQ����\�e��0��L�~ӞBK5���?��>]Y���7h?��	q��&Z��v��0��p�̥A7��%1q�S�&J$, A�*�4����$�2����� ��H�4�U��4!%�%�/DA��ȕ���1��̯*\_�����D���Rjj^J��f��v��Z������� ����K�kw�
«��9i����v wk���R	Na����4�b�>�ªGX�H�����3��=|�%�24.�_7٘N�:Z��MI�-s��f�"Gf�(,�ԙ���\[
�p=��y� �Z	QJ�$1�L�dn��A�!�4�_�diىU@�Tn�Iip�j5�u�e��dj+��9wVh��;I�3�R�k��N�41ά���?��=��G!C
��i�CR$e, G�{�R��k��8��aJ��f���w�E,�m�x�"�����bWii]�?\�k;�}��u}���x.�}i�)�GH��A���9F�a��FK�Z�c੬4��!�.�( �!�n�2& &E;Wڨb�Q3b�AJ3���%Sfy)��"+̳�b�È��I��h����t�Y��ܬ��g&���~1�z�I�/��4i�i�N�6��VX86$]	�O��H���sI�ORxy����/:O)�.I��Et{��ܩ������S�t�.B,����T���:>��%�s���,+p5s}CE�W}��i������F�&��tL;H�,��,a�'�z�YFQ�
"1x�4Kɳ.���|[.�R�0�Qפ���cs���*|�E
�*Rs��/��(Cz�U�*�"7����4��N�}�Y�V�~SHCAf�~��e͕v"���Z�����"�}<�	��L�Z�A`�6J-e�F̾���J�U�WKQ�Es��v(��d8"�s|���=\�}Ra�z�o�������R
}�J pd	M3���(�6 $,�t�.$϶�(��7o�@T!�}\����`�8}Ҟ��,6�1�8I�k�l�\r|'���r��鮿���eT2���jl�d[>}K�-�Ců��:I�}��7��R�im "%�;[�0H��'(�'/���vNc,�0�����a�qL�IL�DhA%�ɖ5��ڗy/M�	���j�tp\���Q.m�I���0���B?��F�<$]�?����ib��֠¬U~U�U̞m�Z�B�^%���	��M�*2�*�8�e����\ifB!��	�L�a9d�}Ȓ�T
���)
��G^dh��E1I����h�4���m� ��h������<����[Y[N�>����t�wϜ���+�v:d" /����ø~�0����I*�O/U\[�q��-N_Z���6QR�;3�=j�
�04�A�mx���w	k.i��$���Zj]8dY�R�#F��<�IӔ8�̖*��r�J�4�Hӌ4�M�=�iu��Z�ԹyΜ�����98~�:@Pi�V�� xp�h�����F̅��9}���ٴ��,�Iӌ$����8IMz��-L���*e�ҟ��{y^���^K�4��y9�E_+�;ύZ�mv���=��.+ko�8�K���͓Yڈ(�*~}���8��1��(~m��6�_%h�Ԇ������;�x��󜿺H�!��j)63�̀7NS��<��i�=���0��UC���yD�l��q�diJ%d���ڭuz������Մn/"���6�n\gei�N�Ǎ[�y����~����7x��w�H+�ûiL�9}���.��0ncј#��� ��ҵu��������9u�<kk��IJ7�ho����L��!�R�l�^�T�*��j��04p����.[a��u��*��C�����6@`�4�L)�4'�S�(�#٣? ��۷y�����[�^�������yV�
�ר7�Asb7��!��nc� �V�8�9�Y�+�V��k'x���\��NC<�S:��N�G/��%=�,Ks\I��D����	C���5���J� ���&�C�����g��ǎ��C>��������}>��#�p��a�6�ܷ�];�3>1A!|��9�vm����A��`���3��q��Ax�Qy�	>����c�l��fߞ]:��#�s�)�s�}G9z���M�:�v��4Oɭ��������V���k A�I�Q(�J�����?���0KGa\�Ql�q���u��Q֥�푤)q�������d�"+4Z���i��EH�\;(�)tN*R
���ڝY���S�ڠ��$%Ir����`���9x�C^}_}�!� �2��������G��o��ϱ}v�\�W����y<�̢�q�bWNo�s�wN���5�)�[��`t�����9���RHO�W=�^J�m�(O�E��DH8|��8��p���*����?�����q�hC��5g���^U��o���^�5۹��O?�?�S��?�)._�Ɨ��m~�7�����:]S��V��������!�j�
B"� 0����u��p�l�!������ n�Iu���&�S�4�V��"�|N�����}�}{�����_䱇���������]~�w��­uT�����v��Z	���u����{���W�<3�&QJ��t�7�o�o�}��3�s�:~�K_�7~�+���Y�`h�����#9�o;��s��s��Y�(�6��bs�?uy٭#Ah��*�J�+���������8}����J.C�X�Yk{�<����v��y������0@�4��xe�s������SX�PJ��*JG�Pv���v��_���"��G_���+d�ٙ�yA�$LOp���|��g���&N"��S��^Q}0�Fټ:��H�:�����&׮����W����Z�R��m���0@��V��m�<�ă���}��{w��)�gB�����r��[�5~�����_;A�2��YYn�H�}�v����O|
]��mD
aȈ����ƗR��{cݗƧ�|��7�_�����yk�n5�$:�B��&3��Q�h��n����S��43 +r�<5�86�xˤ��QI�D��]@�
N_��?�_�����^�y'��9�G�y�������������˔gs��ܘM+����_�Q�������+����>�fwt'ʖ�l�o�~�O13=Al� q,�����/�����P2ep$$�$.#��y�1{�A|i�Q��L��"K��4����5Ef�q)%�硔B�9�0������|���U�כ�hk"gR�D�)�&�;�L����=���x����'��?�q��KsǺD�<�Iy�.8s�
��_����WX\^��̻P��3�<����Ϳ��ٹ퇇r�����zq���[������p���06�{p�B|����ԫ�5|��ZC9H�W�l|`�[�.��N-~ m�D�.�#�R��ن(
�u����f�{�C�L_�R1�q��J����r�&Ib�<�:k<�%I���z3�S�A�Xt�����8���I���� ]�,/�c�aɗb�?�s��ܣ9l�;˫�|�������5ʌ�f��۷��c1::L��1����6>1k� ���vM"B����x���s�,q�����;�
�d�����<�7ϭ��z��%�1�VHaq�ZaL�3��P�|'�s�erC%$���q�<DJ�u��&QJx�3�,�R1���:`$|�'�K���S�5����d�T���z���P��]�{��J� ֭�HI�4k뭾3�����4��lຒ<K�M�%N+�Ҡ�������ѵ�������������:��`�g�*��!Jk��v�+iU�<i��w� �<!�*~!$Q֣ӊH��x����m�֞����LCW*f�T�j�� M�n�ւ��	��1I�yn<Y�Z!�^|�3�-3�̌;�����N,EXGI���o�i����B��F�Ҋ�@��AjH\zQ����{t��˫�I�w0�Ω,+����!7��cH��('�s*u�7�稛Rd�j�G+M���v#�<�q��1�[��3��K�}�Z�.c#��ۻ��dblԸ��y:�t�U�*R<�!Di�;�^��w�r��-�V��[~��"�����&�2��:ƍ���HA���-b��
TI��gd)�3� �ܖ�,�\y��	��O����]��Y��:�#���0�m��g<~i���6��û���d���q]:�.I�048��F���/s��-�7�H)hw�h��������5E�V7�h�L�2��D�%fItCI�d,.���oq��ez��0��*F[�g�g�o�$IA�c�y�O����L��:��(@��D9BhmJBIa�׿�����/��}�y�WV�תw\/��X��Vx��w���BQJ�yfo')i�Q�U)��׋��)��N�l��	�mT�V��e9q�R����ۋp��jz�3�<��!�MO�}v��;f�~�7n�frb�V�ˉ��y�7�<�7���c#�ٟ�1>���8�a`�����BR��)aKp���'	׮����+��7_���K����n)}\=[����266��>��s��G?�a���fÊ�<+(,1�16�B����݄C%��zۦ��%��������f��q���(�w��{�#�04�$�;��$.Bo.�[�=����*Q���������"��DqJ���)��,{��7\ץ(r{m����@)�stB[d���Y���*'�^d}����o�<���F%(-�HΜ9����8�ϣ�g����'?����[������\�lnb*73=�L5,��p]���&��a���������1vw���F��
����O}��>��f���U�^��֭[�z�]��P�0RH�GFطw�g�)����%���o�����������(G���ޝ�+!hw{��p��/�p�m���>�����m�3J+\��Jv�ZA+S��L��I��B�86v�Oq�����.��~���l��ۋؽs���GXmopca���I\鱴��k��F������O=˧?�;��Q��/]�ҵ묬��h��
%�O 4�*p\��`��3욝�R�p��E~�7��o>�2g/\�u��t��a�5S���~�O|�i����uX^i��/���N�:IVh�-@�;%NRv�M�>�g>���݅֊�|�u~�w��/�[h	?�����]��ǉ�	<�=����9��]��_���A�5�����ǒ,6F۽Ę 
�4�z��h��� �z�f�J�HYQ�e=ҴC�:l�Sn/,�jwɲ��ɟF�<g��`��<p�{voG��7�:�?�2Zk��0��~��;��� yV�ҫo�����}�,�+��*��j1���(t���x���̟��c�TB�\�ί����_�KKk$�ٙ�U�*�̉zC���� ?��≇��9g/��_���_��wϲ�֦�1��n�G�}^�v�����4�Q� t�����ɇ�s��2�~�e�|�-Ξ����K���0�lp��u�$�svkaY��l��P:C;)C�v�Lr��~�?��cvpd�v�a��4۷M0;5ƶ�Q��ٱm��m�l�evj����* \�� ��2��3�RdYf#x� �fj|���m��f��9>���|��'bii�?��s�����w^|�7hwz���=ڸۋhuz,-������F����'�$-�.7o.��tq]�:4�KB
��@E��216̃��x�F�N���_�&��ů���v�0�!�c��~��K�ܸ�DG�˾=;��SN_��Қ��ԩ|�;/������7�8�o'#�ߺI��ۂ�}��RJu��z��X�};�q��n�=��=;صm�٩&F�l2ج3ج2<�`th���!F���6�69��� #�|�-UE�FX�������N�Z��>�F���!&&F�٨�I�ع��ʭ�e��ɣ�ȡ}$Q���x���_��y�ť����ݾ�T�EQ���΍�K���mj�ёa4���uN�:��ںq�W�fIJA����%4j.�gFx�чh6�>{������ݗ^��Ԍ�+���~a�=�q��p4�<�0��o.��ۧI�����dY���{���adx��GP�֘�z���6Q�n���f�71>¡}{x�y��a��c�Y%�$
M^h��4�r�w��ĖF��u��dth���	f�1<�%Z�Y!MX������3ӓ<���|���>���$R�,/�s��<o�{�k�o2;3��{سs�KW��o�����*���kU�G��/��q�: QĽ�����D�u.�;˛�cm���H<�,U���R:Hi��bm}���5ڝ�u܍���=�za��4�ۍ)
�r��*Q��n322���s��>�;z�G<��`�8��v"�Ԧu�%Zk�4�V��w�v9~��8��=;���Q�d�5`
mH�����$5޼43��րa�p��h�sf���������u�;�5�/4�'��$�FH�Rm2p;������-��F�6F�1k�Ƶ�������b��)�V�����H@��,k�Ja�$iJ���x^!c���t�2��j6�wܔ�iTHa��=	Je��mn--⺒�3�4k4�69��fcu�������KM�U\G0�m�'>�3��s�4}P��d��C�SnX��밾˓WK��^ܥ�p�˶�9}�I>��s`�.F�ǽD
Iu�y�*o��.���6��_���A�I�Gk��	���G����8�{FmQ$�	t�R	C��7!qZ��#�����EA�x�K�n[�<&��h]��������-n�,���3+R�,ꯑJ%&QBxl�l��[����^��ų��֛���}���6��+���MosQ��:�G���G�8����cd���&�Eil�Z�I�Ph��W���4�U��	��$I���h�	��z�F5�Ъ��k㪄��>��y�������uM&j)�¾�Wۼ��9�����[Ͽ���2c#<��q��S?͏}���߻�Z�bR�,���+�zl�J����D�{
|�?y%��c$�DA��&*$�)q��� )%/
�"5�U���Q*�����%N��D�����������QBШ׶x���TJS�U�1;ͣ�ء�L��HI�
լ01z���R�V�74�Mfdd�����&�M��h6:,-/���B��	�*PyBՓ��>��#{���n�F����r�<���(�&'���Y���^/fy��F�>��0����p7�$�ƓNjw6x�)F�y���P�u*a@�e�q�eT���w��]�4ԤJ� �8H����@H�F����8��0dnv'Sc�
�
��5�M���faU��3<��q�>���(�-0j�u�,��9�Z���f��b``���a�����l�WC�����u^{�u^y�U�W�G�VC8nl9=1�3����ZC��,�ٹ}�?���������޿�ťU~��������o�o�s�v�l�\���S4i|�oZ\���)�,l�����qb��ww��T���i��fﮤɭ�6#ϫ�n�$hxS7���;���3K��	;�s��051����x���8r`��;�SO=α���FѷA�� �$��U�����]�+ʲmJ�t;�a���4��ӌ��R���g�����T*�&�����������[���[\�t�^��t<���=�e|t������-ٳF{n�ۜ�t�W�z�S�����@���	��Ů��hUp���%��s�*�^Ab��Q�hE�K������|3v��]�UdyA�Q��)��1ѱ{�XH� m���)L�l��/l�H�RB�4�Gi�ERv���P�mۦy�G�97K�8�z=z�)-���Y��w���031��7�r��E=��&�v�bff���AkD��	�nnᤔ�j5F�G%pC��.�����;����\�r�n�cB�Z�H�a��mݿ���\�d�:����/��_��7�����[���|�ɇy��cLO����=��]�]ǥ�TiVjT��l��4��6*ԫ��ſ��0o�x�A�
!(��4i��'i��I�!M�V��||���{.�,�qU_�¹I��K{(e҇/4Ν[�s��o.������K\����K�o�dai�,˩U+�����8G�glt�B)�B!���W�p��e���&&m�$v��%���<j�^�Qo�طw/�SS(�X�u���z���6'O�bcc�T��4˨T���w'�Z�NIl?/<VVb�}�4�N��ƭ�Q�D�� ]h�,�h��v.��㺌�ȱ|�|�����'�:�ǟ>�Ǟ<ĳ��c���6��J1(���b�;#J$�vG�� �V�� �����wΰo�8�wO�o�6�����	�f��팏�#, �T�2��\uZ^Y��W^�ŗ_����˷��.�=�o���Wo���Mc�<��涍�kn�Z%�����(��,ϨT*�l�ap`��fTv��|)%y��>�������:t�F�IQ�DqL��dJ&EI)�4lrp�cC)�f�����iv�ΰ{�v����Ԅ�)Ԍ�940����A/�wf�])�`����O�{�4���1;�ιIv�M�{�;�O06\ŗ¢z�͜MsCLYJ���X��2���������!��!�*����x��Ny��<t�����S��Ï��dn�^��K腶��������Z}�]����y�����s�}�o?�n_�M���\�4ej���a�B�H�)�<#�#�F�ؿo?���^��m"����EYl_��DQ����9�x�	>��Or����fzf;a}�|˞8�s*�˞���g�� �3<�gnj�����G����4O>r���!�MFG	C]¹�@����G�""������J�J�JV�Vjԫj�:ՊK��q���G�+C�5}�_��0������1�YI��8���Z������h���	�F�fx`���F��lzT���H	l*S�QǑ�w�exb���Ó�O�2<9���$���4�ukR���1�M������eQ������$�#���!J���]+U~iԕ�u��l�9fgg��G>�ٟ����ȟ�����O�sn�IC>�Q�h`vz��3C4����7��o>�
�.\�w=��_����c�~�]�V֨U*��5��
AP�U�UB�F�ɜ2@�M��A5=F�}�F<Ɔ]���}&��n�n��Tj�
��Ш�h�)���H*t]� ��-n�Z`iy����<��Q��8^@��1PhVhTh�4�4������`ͥJ4�n��K�z1�o/���h��9r��<ƃ����#<���<����ڽ�F�nӅ4�f���1���(��>�!*&''�>����1��Ͳ;:��h��x�����K��J�����y���x���y��q�������j��8�8	�2>6���1[e+a}�Ej9����`aq�$��EN�e��6�VV7XX\fqi�N�'��>ҫP��4P�	�U�f��@�c���0�P��8�Yom������"���q��gvj6,��9Ea��J8H�\��ko�����:kĽW��ع��a�UEj�P��J�PP�jtZ=.�_��M��
�J����x��wy�����C�=���سc;3�욛e����������Wޠ��mv���bz|����� MS���±��4M�3xkǗ��߭��%����'I�_�� K����9.����Ԏ9y��z�g�y���SLM����'���<��#>��v����z���uzݘN���'���gYZ^�P��|-�����L�ynF�i
U���������۫\�_&�
(��y��;���\��H� f?�W�o�)7o.q��e.]����*i��
��
��;��3�TC��&�^�~�u|_������۴�I����̙s�9i�ۋ�[纬m�Y]�  �
����_���S��t�&��2;=���2k��{n6��Uvn�We'n��[��ݚ���|)k�m=g9آ^����W�(��v�ͅ��hr`��<��k�:�^��7n.r��e.^�F��cu�ť��8w�
7��E�V��Fݳ��� �)�GU����Ÿ.����5�\X�Ŭo��|�:g�]���ڝ�|B�s����M�t��7n����9B����@���#;��nzy!P
�a�#+h8n�rk��WViu:�.�������V��i��e�]�ʵ���^s��5�~�Ξ9K/�4��NOr`��Z?�]JI%����K�\��vp����J�:0���[��Rs�� �"���8��m�:#�t�r}��C��O����k��p�wN���՛�qF�d���s��<��k�Y�����sh��A��G�H��8�Fz���ҵ5N��E����ƹW���F����9�Oz�H)�VB*a`�D[�G�o�z�R�BI�����6E�L�-����3ӡZ-�ih��I!�h����y!�F�Z�V��n��N������CV��j�J�b��eG�̖N�{旟}��r�o�����u�����l��q=j���*K��<���9s�*�x���NL�iŬ�nб	+Br�j�B����-���ߣ.1PYb���Pu��ױ����Fm���Z՜��q����w���H[�^iA����"t#��.��G�&Y��D����Q��FssN�o�-aP0�Lϕ��@	I���=�%�}C:d�����١�G���S���������ڰp8��x�K��,��G)�����8�j�"�,wh#K����ݢ�$8��M�0�h66��N��a�j�����!�۠�\�d���"*�T֨�mW�Zk�'PJ��$�eҲ��R�V� UddY�w>8� } ����B��&���nڬ䱳�����׽�l����[?3���\����������s]�u�Mwϲ��ȑ��l�\��:[��?@Q8�y��|��@kAQ_01��WM�o�{��MHRž�ٷt����6u���*�F������	��#�z�6������y��M�q���6��s6hXI>��)��s�DI>��3�.;����#���*���� ʤK�u&�e������$%���M������j�h4�TB��u (-�4�%���TH�p�����i=A�c2�F�jP��\�4��xG�����$�<t�a�x�~��@�N��bEBh|_#�0�������V-C����������Gx��xྃnj���LV[E�I@T�g_��3ѸtKb3��O*��n�n)�YEf�u��$H�1�f9y�����Ȋ¸x�L�rЏ�48�o;O>r?ǎ�g|b�19�����e�֊n�KCz�G/$� /�@RBg4j���#�<ʣc��$��Y�A� S�UQ���g������_��_�g?��l��F�$DqB�k��="g�ԟ3�:a��;�0Y5q��عk��������?��c�9��o\��8�t+PEB���[j�9�!.Δ���T�w�Px�5�-3x���F�ߓ�^M�Yg1Jֽ��]��,�`ʝ�OO�&�d�Q������,����E���	x�(������P(��VS,t��_a~e��KMn/V֡�H4����61�'?����5��/|�'|������rA����z�o�N��ˮ�۩UM~��:8�*�xDy��v��V���`�[!Na\���P�j-dߞ��ݽ�]�gi�MEdaH�8&Jb�8#�M}_a�@�t�&Ź�)e^^���nm�j�����IbJ~�Ê������F�9I��v�t:t�]z�I��q��3�ȩTY�!+4qRKۦ�;R΁ ���daB&B��۾�����k� �@V�#M���2#Q=��]�2�VV�Vn�UXZwY[�YZ��JHs�*�c�޵��;��s�~��&�a"�c3������t0�ܫ�����<�h�n�pme�k+\[��z��� I�,SE!���̅���;�%y��fII\@�m�����0���]D���U����;��]�^�ܲfl�X�t�=?��9�cz]Sr����_�N��ף��Y���#$�q�3A'2Y���T(��T��G�wh�]JpS'^	dQR�ZM#
R�c}c���:��V+a��Y�VY�lld�^��ʈT��E)�іg�����"�0�i�&��L�b<�JҔ(�$�XY[cay�յ��՜����.kK�+)�nuX\�5j���8`���yV���&|v�M33=��� �jH��>y@��v���-c!L��4�_��9����>@�-����}��<���zlt:�ij�r�|V�{]Zk+dI�k���ѡ��XY����t{=6Z�#���µ�Y\���hV�۴�7�t{�q��2(t�m�b�pD��3̕��x�᭳��&}�}����o��` Y�M��AQdyүr�u����!N�(&K5i�IRE�*R�w��э���9J5�Q���\&'F9~� �?|��c���o���fn�6GE1�v���:Q�õ�aAE^��F��E)�4%�"���9m=rqǱ1Ƭkv}c�յ���("�"�^�<3c���no��t�V���l��Ƒ��ٽk;~�36:��y��1����@��c\a���7f�х$K4�NdRk���uZ묷[��[�m���h�ı�|���l��>~x��aU6�Vr��8����{$��5����lXi��� !����9�B����s�>����4�<��|�cO��#�	,��у{��'��Cz���	�(fqe����5�L�A@��,�����D��%EQ?�Rv�VU_m��@�lц��EΜ;É�'�t�"����|w������mn]a��������3��~������{�,�����G�K���g>���sT��yDmI�ŶY�N�V����9w�*�/�s���]���KW9ui�ӗ�r��V���/�X��3�A�wX�.lQ���qq<�n�0{m�fH)(TA/�X^[���2��z�:�W�rm~���7�zk��7X\Z�׋�8T�j�q'~<59Ɓ};Y\^���|���~����o��F�=�g�65A���F\�_���[�d��˯s���~�-����l��$IH���[:M��N�r�?��{����<�<���7y���X\^4$ξ�����f}c��7����R059ƞ�;(�.�/���ً�:w���r��%�_�EŖ�T��R��$���
����y��-�>w�wO_�w.��[�x��mn,n��fy��\�r�Q�F�Ԑ;�H�I��	���` J���ʹ+79q�
��]�̹+�<s���.s��5Μ�Ƶ�K��BR�,��}���&#Ã\�v�/}�;<��k<��+|���s��"C���#4�U�8��U.ͯ�����Rx�G�Z������kܺ}�$5I�h�k�iԕ�eYH���ĩӧ��������p�.^dqy�$M�o�v��f9�n����e��"��4�ujՐ˗/���K����^z���*������,-���T���xGJ�Bs{������X��Wo��vs��ז�rm���-V[�n�a, �ɦU�)R:��I�a6�w݉Ƹ%���X����|���}�&'.����[�q�:'N]�͓׹|m�!�)���RG�Kj��J��)���k��
�F��Q�]˲��|Ӂ�+�\�r�Sogɓ�)EQШ�ٻgS�S��������ӝ�lU[�+����gϝ�ҥ�t�$�#c�?p��{��mr�1pf	�V7�����\\����,MY[Y�������%N�{��'Np���x�].^����z_3}�a��q`�qL�G��H�j�1�>��h�{<f_dɶ���7H�cx��\u���'9�^J����t��^R��e�:1�('�������R��.I���j���mz�g�x���ws��^�x�~��F̺��B/��}�괰���'�ska�
|׷����1=��z�n-\A�^�Z��8&�,���K	|���&&'&�9QbhR�'�8p� ��w�3�T*վm�:�5���s��56�=S��q�t:�^X$B�MM099���33���mcdd��z?�+,�v/��֗�Ҷt�ua�����ջ�Fz�z�R�g*>h�H)|�F�Jxx�C�R	}<סZ18>!�u<B/�;���8�XX\e��"�##|�Ï��c�y��x�hֹ��¥��h�:T0�t��>s�s.���bR�\�4�+UFG��6���%f������t�[v`��=>���8�cC6f���;~�C248��Q�ҧ>��Μ�����if�Ď�ӋXouصc�=� O=� ���|�#���=�C���؈aݲ�yw���{}�)F�����@�q�'��-ȋ�4mY��~������b��S�gi�eQ�s&Ժ���׾�</��:k={�8=p�4�x�W��7�K%��Iu�����W�y�����9�4���lV�;>C�4eqq�˗/s��Z��^�'c�l�Lu�8���h��R&�'8~�~>���<��#�݉�yDqL'T�*����^���\���[�±V�R�z��ܶIv�M��x�~�A9~�G<ƃ�����T������BO�������J��Nh�������2S+GaS��!@z6K�}e�[�2�'��Y��:��uRg�~)���TQp��o����K�X�h�g ��eQ�z=���XYYacc���5��֌���!�cz��v����
ׯ_gyy�F����{9v�ۦ�Q�T� <4E�q��o�����7YXn��p�֊Z�����(feu��o3UF%p�%�}�,G�Z��q���G�<�>s���G�YC�J�lK'��H�U�T)n��U�L���Q�p<�|����݀�WE���e��CO>�G�~��3���;���I���У<���	�o��Ĺ��
Y�r������x��e�<õ���<G�͆VJ�j�XZZ����,..���d^��,�Z����\�r��n����A���I��v�MQT+��ga�6o��/��K�+���%a��'�ï~�W_}�wO����y��9{�Y���}�4{7���i��,p��-���y���g?�GdQ�V�F�R)E�9V�L�D��[��0�ŵ�q��jB�3��rl2[�]S#����m׫,77?<����ݴ:]������W���������^�����#��g�>li�u���������ۯ�ɭ�%SL��޲w���`fP���6��u�������f�lA��*��O�s��M���	�:y�յ���식�iQ�J�����ֹ~c�k7n���b��%M;Hi��Z��n���d�yVE	�^lڴ�����$���¢�{���%Cʬ�Z�L�����C�2�@�] �r���	�I� � )<������s<�\������l�\���Q��B�if�ql�����
���8u�<�<��/����:�*C�*��,���@5��-N��ȷ_~�g.p{q�^diN�8����T�B]"rU�F�{�XL�I�0��V���K�y�3���Y�\_2�|W�^��F��W�}���A  �3�^)C
%Xo����u)�_�c�g�o�Z<���$A��

�yo{{���H��Y�=
ep�,Flp����\��� %����}�A�66Z\�~�Nw��ah6���R���I�V�45��F���&C�M��f��<���T+!��n�ֻg�҂�������*SSS���0Ьs��A��v�=�G�F�[� �3�ֹ��N7�q]�U*�O���o��l��"c-\ʱ,پ��%�5��^���y���I�_�j1�!y/�*��
F�����b�Q�Q3����tㄛ������w�Nv옣��x{��V�dr���x�j���p��	��Q������Ԙ��3<�`pp�}��8rp����p��e^~�mV�֍�ft��q$N` í��=���#���W~��m�,-����or��<E��ē��&+%Y�!�͖��u�6=�Ǟ}���y��i������\X�G?���7�:�0f[Oۑ��)��K_�&�._�&wv|)�B� j�
��욛`����S�6M�c����(k�!LFL���!4ʳ�n��z�7ory��-���N�$}��{��$�w��������4&M2�062̵[79q�,����z�O<�Qq��9Μ��z���J|ϸX�<�@���l��2�Ab�@r�m�ڷ��v3�&_�ڷ����W�t�:C��MfK��Ջb���}���W��3�[Ȁ#di��*� ��B����=D�d\�r����-g/^�cO=���0�w��)|�o�����-n�ZB}@��!Y�%	�j���Avnfnv����I-t�T�x%jW�4��Ρۍh����r����\�t�V�so��{�R�������?�	:�k�$��ێ��у�X]_�S����>C��ձ�-pL&�V��M�i��1�	
��_�Յ+���s/��~�7�pi��
��"gfz�'�����>�����Q��_�q$����ZJ���8&Ҥ�]�M�iKk��p�^�z����_��F���TB3���f�v���5��Ґo�w����XQ(�"�q\|����z���AՀZ-�Z7N�r�H�n'�P�(�Y^Y"Nr�B�nw���,��]�����R�4���ӏ�#�x�_y�w�=I�Y���P�5x��O�`}�M�V����|���h6�ifx��1J�5M�	iʪ�T'�#M�\���-]�-� \�4�w^|�_��/�Z	�[�`p���s|�Ï1=1F����^|���̰t]ǖ��x�c�TM��HJiN�$)��|㹗y��Z����#m[�q��:�'%Ȗإ� �!3.E8	\���^d��g���,��F��L���4����c�'����[T���8Iy��c<��ü{�"o����G=�'&�ا>���0���$i���0?H��뚢�ya�礀�0�G�	�]�1 N��!�d��u��^\�������,-���޽������`����`4�:�����o4\]o�iÍ����Zi�����5YOR��P�WUHG�vTn�~�h��+�
& ������,��e��,3���J��vD��55�=��,��v�˾=��Гq��^ڭ_�����v��������׾�<W�o�e�C6��_���v��f ���HSK�|��Wek����So���m�������x���oo������'Q�Hʠ��k����&���<y�u��EaR����sld��r�+5�U�~�5��'245vn��3O<���(��k�O�����/��}���6�f�n����]�o���K�v�+�����P��O�_,bˣl9z�1���������n�r m�l���������� ��~�5��'S�SJ�Cvq��vZ����捷O���\�v���L�?3Ҷ��<��|��$wj����_I�^���PT��LI��}���))5nU��"����p�"�=r-�������פ=��U/'���yϲ��D-k�f=I����d����������<IҾ/�O"w��?�����u�?�1Qf��k�m6�������u$�e�����Q�:'/be��EQ��n�qS`sK.��C��j�AhI�l6��89�TD�Ga;���� ��)�|�R8��G	��V�Q	�|�y�(\O@�#0еn/B)E%�up�Պ	F٥n뽛�09yn��L%
�x���k�2M�X�������{��O{�֗K��B���G6.n���қ�n'�*d����e�wZ��h[��n����J+�� �I���]��*�n�萹���]�1���z�R�)�ZO��6K�~�|a���.赔%50תV�>�ltx�����}�c_��I��3L�ږw/(J�i�-�oK;{���O��'����H����Eb���+Ra�D�4�L�a!5y�IkZ�Z���a�,a�բ݊P��Z�>3���0N��Zo����ʊ��y��t����f�z���`��A���:�.�n�du�E帮����wn�ҨЍz\�|���6*7��&)4��4C�RJ1;3���#Ct����Yk��H��Z�յ6�m�tS�ݔ>�261�+\���n_���PdF�:6=�l{�@3��XXl��!�0�=kUV�7PJ�lԙ��f`�A�q���K����0����G�����M�7�$��Ǘ����6<�KB��c:P+L��kt!Ѕ�f HW�2sLX[:�wV��y��	>���7�FK��x����3ڷ�=�瘜ax�I��hw�b��V� m��EQ ����8rx�fdp�J�Sm�$IJ��c|l����sp�^f��s!�r:mq-2V��Zc��#}����ÃTkU�$b��8z�a�ִ�B�ett���I�*�3S�0��4jU*U�5�nd�i3
[s��<��Np��Z݈��6R�f�ٻ{;E�hr`�Nv�fzz�ɑ1t�cf�M�w�����������t��"��f�ڞN�k��y�62�K�
Tf�K����9VW*j^
��5�;�taʅ��]AQ��w� �/�4�&'hm�8}�2���Ǟfff��H�q�*�S>����V�7h�� ���sE1�R<��q�ۉ/V�6��Ç/pY^_�CO<̑��r���:���Jr�ҼqnX_���4͘���C~�#�w�Iɩ���Ӝz�A��������O��*X][!t3��Lrp�~j�:�C�L����A�e<���45�o^'M2Ta�馽�Mrp��y�1V[-W�q��у{y���T*Uf�Mq��.:�U�*BJ�5}��&Ƹ}k�$�)�n'�ۉ�`���6K�����D����������������dԬ/)!WUH�����$A��*���3�S�۳�ёa�(ac�͵��ٱ}�<t�[��x��Ӝ={�0�0::���n/�ƭ� ����R{�C�M�\���o����"���R		}���B���^}�3�/�b�ۅ�8,���jw�E1B��@�� �8tp7�=tk+�{�<��_aee�^{�N/f��G����jP����ccf�kȳ�w�~�kW�9�o/a5�G�Z=z��X�%��bjb����n���1����HK Y9'�=�ɓ�XZ��g'baa����"���h�XYݠ��dY�1����ޢ��Z��Kՠ��aL�Q
�B�+�>%���fH�ɔq�
;��j�?� ۦ&8�*���ۋ"��f����{����{�����0�Uۦ'HҔ��.!����{Q����ݏ�7O��_���Uf�昜�`��4�C.^���}�;̟�L/�ص}�JH�7n-���A%4��B+�G=���{��ݗ��;/�F�w׉:k7�|��n��Ph\ܰ�v$yZ�	˫����9�,�s�S�׸q}���~�?U�//S�U�����n��h4j����J�$������;�9q��[K��O`'��7���o�[�k�������v������"��ھ���n%�0uSzѝ$�aP�2`�JC�{$��vma��B�s3��5�������Ͱs�vu�N�8�L�a�#�$!%�=��i/��� ��)a�#��f_^i��fdh !C��k؂C�8!�s��H�{-�A`�9�8Wt��s���~>��O�3��i�;r4��0υ+�IӌC�v1=6F���fK�:f�ı!r��h������jU�Z��nK���˞����܆vrnݞ'�S�,giy�8���`ٻ��z:�Jx(m�|MZW���8957E��lJ��-]����l��n9�g�+M�"��й�kX1�����1Ь�NP*��=���l�Qy��� �S�T�G���ނ;��ym �si�댌�3>5���(y^p��"���Rk01>J86��� �BH:�Yf�x�R�8�C��yQ02<�����0>1��c�صc�f�F'N�p��o.0;3���)*��=8�$�Vh24>����㰶�A�df}/'���*�(���y�];f9vxB��3X]k!�Qi4#�(�V�0:>���(�#�5i4�������ĩ�����j%��<��3Ǫol���,|*��S�,�J��:l�;x�ö�q��(��o�N�!�G軄�)��U\ףՍ8��Q�=���x��yV��mꯋ����2�����Ћ5��L�l�c�>����{�MFFG��jt;]�Ր�m�<��1�$��w�p{a�;!Jآ��ѡA���N�Z%�
N�:GX	ٶmʀ8=8���	��V��G�b�٠�j�)J@�iE=����'?
Z��kos{a��F��vt,�u�����=�� �g�y��3|���gtd�];�سg;�˫t������� �#ٱc;�z���FGG���*�#CS��BK2����w����v�$��*�����<�01�2c�[�uxh���I�U�+W.��w_����8��6Z��\�Ѩ1=9���Sct�=^}��n��l/%����n�f�M0<4���c#C4t{o�u���=CQ�����v�09>L��8s�'�\�Ƕ�Z��}�Y�F������LN��#�|�:��+y�ٳ�X[�23=N��cqy���U)�1;����CC�qƉ��9q��ȡ��j�
yaB�ӓc�j66ڼ��IN����H|�c�٠Q��}f�=����"._���:�kf�'ؽ}�f��z{�V�Cm���ϒ2k}�t���*r�@aǄ�W� �mz��@����;ݺQA؛����̙s�9u�*k]�$Ei�ͅe._���4j4�h�9}�g�_����&D*���]3�q�
)��8y����wL�caq�V����q�,�䩓�<{�ť�xަOl�҄�5�l6 S������,�^ �;ܺ�B�����+,.���3ԨS	�$���Oq��y�W�P��})RJ��G�3��.�v��W�q����Ȕ4-4�*�Ãh�ҕ�:s�^��w]�ML�n��7o���!K7��XH��i��6�91��q�8���"�reU��f�Wjӥy�� �(.
c�a@�Z!I��Vf=�[�EQ�%#��Dq��4�,wE�H��1u�J�d`󼳼 NL���[߽Z��U���Mr^�a���g��'�sk�V�TB�,�ӋH���#m�кF�=z��똭���`���~���5q�w�����-)�0�Q���8�Ӎ�c���ת4�[)#�M�έ�W(���D1��q�HI 3�+<�6����ʡ�+U���c���*�Hm����81��j��`٣8FY{�"�=��b ���umxҀ "��u\�8&M3�6�S��A`�g%IJ��i�����Sk4�|�;%/
�����x�����>�*� GJ����� �T�#��?��n�ve|���M����>q���2H��s�4˟�^Y�?!��IC�wW�ޒ����=�Ǘ�2��ff�\�f���@�i؋�C+����B�����sGg�rGǗZ0�O'h���s�-���p��3����uSEr�x��k��O�ĕI�keB�S�W�pq#��Q��0Q*GI���h�|�0�C���F	�#�aw�9�=��{R[��2(������r�R�
�J��*�m<���V8�'i���=�0�V�yf�&PEf��B�I�"+��:�T��\C�f�:{�?~���,mPd�ZJt5Ef�n[?��㭔uI�(&��50�ɑ�i�S��������u�&GAlZ��]�5��)�iD_�Zv�*P�G���Z�H��&���=\�6�>Z���n��
a"���JJ�� y�FI阸�e���=yB"��O%$Z�����O���2o^���٤=��)t����!х���=����� �w���:�A�o��Gv�H
E�Kx�{/����p��5�^�ϑ3?���+����=��.�o���U��b5���MI��d)A���~�Y���7�<+�BjG�`��w BE�GMH��6��PK���c���^��	6���C��[��w�=O
�kp�}�R�-�)@���Y>��)�g���8W.L�9`S�@����6T2�z�e����s�,�v�j��k!֥�=w���3��M&l�Hta,z"�<:&��n�\>�#���������1��Wy���XZޠ($ʒ �BPضz��O�5!��p,������%����$�LP�e�&�`ӳW7�GH��
�*s!���l�0��@��Q�噻s�B+��U7�F����Z�y�D��>���d;�B�<Z�|	{�M)��B׷�9..Cr���w�o�v�<�[/��?�����/����}Ϡp��1R����-M������ī�~�5aY�_+�Z�r9��O�q��Ï}�����162�;�N�/�ݿ���+���̅E�J��4B�y�Ҷ��9v��� �������"���%{�O))Q�0�@E캦Åij�@U3�p
��}#���}#LA?����|���8�j� %P��b,F��?�������h���#���}F�����)4��������9s���^�� j��3�f~_�n]����'��B*�]��1�4�eh9v]�_u��O~���7�*�C����;����_�։�d�	�x�G��`�!��ގT��Ď�:9�]���6ٚ�\��		����@�Py�p<��x��ITa�[����n+�4���%\�Q�����<�w+)���l,%���p�dx<į>Ҭ�{˭6�+���`���	�j}�J\$8�4���DĨ=k蠀\�g���20ul���"׬.ĤI��[�^�ɳ�_��/����ߢY���˯������S�h������8�8h-h�U���#�����/���*J;Ȳ�5���\��FR�KEQ�yN��ۿ�O|�i�:7o-��^���+�lЬ�N698Wa�L�Ω
ۧ���,h�a� �a�H���Q�}i�@#T��"�-蒤��O�L�N:�ǡ9�i������b-Iһ����=�v��[�ꪮ�gh{<x�3ƶ��%$ca$x� ��x�/l���~�^@FB$F��g�ޫ�o-w�Ξ{f��֭��yⓢ*N�9�y32�/���OgU�G�VXe����MF�k���ԭ�!�0n��dA��50XrX�lq�C���_5.(:k�גA�5i���ƪ �`��"��@����AF�<��u��X��zͦ���XDg-:k�`U�u�c�r����ɐ����^����s|6w���?bw��ĩ��6�R�FP�qﴮ��Vg���kfh�EK����%^��i
B�"/k��еj>��𵯢l���!�~��6�D��W���.�WCn]�~a�+���p&d���_��]Z�-�q(jI��aD�')#lW�:��K
+R�Sɥ�+�xq���=g�k>��M��z\���+ԙ`j�ԾA�Qa�ı�՚z=�vj:���h�o����;.�D+
`�"P�`i9d�)�ٴ$M+��p�3��2�������^��5[���r��Y���z%`��1x�<���e���"�K���EJi�y������x�ǣͦ������Vm`���[����|r?��n��7��T(���,��ظA�<xt�Ì4�D��22�4���9G��:�ų<:���G�}�i�/_���5�.�0V����d.����>�>��G�<L.�[^`לe�\$���GW��;m>\'�\�����$�m��U�{��9ǁ��W6����^`�`�aaa	�n���NNbr��<�x=����(�DGfu�*Vυ�6"Z�Ld|���8|����1�N(k���?���`�y��tj@�r ZP�����r��ʕ%����.��`~t o�Qߛ�?��(�.b�%r��d�t����+_EI����|����7z�R�l�=1����V|��o��q�����M���	|��&"��yp��?��[T�%��vp�:pP>�?ネ9[#Mn����!>[q��Y�����1�7\�����E��Xb.�2&<�	�a�5jo��;���a�s�<u���/c{穃��%8.%�y�x4`���h��8`'�aL��T�šC=)�U˪��x ����k�]Vn)2r6����[l�7a��s���ѣ9E)�C�ΪC'lTF�Fr��sc��i]J�S�.�\������R�&�wf���A�{�ܜcmL`/!ql�Zj��d2J��������<R��G���w�?8ni�\d7���[�}+���}�����s�K8N�9�:����,c�u,��3 �2�s��a9]&��ݭ�;[1[ÒR�z"d'�G�O"��a��>S(�
K�x(4��t��(\�o	��O�kj�(��l�9�^�G��Nϡ��E�e�ófI�<����1���b�ar�$b�]Dm��oKt�󬽤X�Y�xtg·2b��!�a�.#+�t���5ڲ�sqz�x^`�|� ]5J�8q��ˆs/G�*����79��v��D��S��&(j��QY8k+��`����]|�Ͼt	%�6��[?fo�������������v��Փ��/��7�(��Q�(
�.^4 �B��|DEm�K�xQ�ĝ	��p����%�"�0D�������
ʔ(��#�����A7�||�����'�x��x�.aGv���!�]:f��
��^��X����Y-9��!Puiq01;,P���^-�^�k��霅�N��;c>�1��+���E��B2�P�5�sXZw�;z*)vm��&���k��i���u?������c��M/�����8���L
��Q�@�Jf�9�/��s׾�o�lo�����e���</�D���]�,�����T�K�����#� r	"�&���i��ߋ:��Ԡߡߋ#� �#�^'`��J�nH��>A�C�	q<7�� �sp\�)}���q\���8����N�O@(zD�G�+B��sl�4XT����\��{sJ%�f�;�8h�`ٌ�u4���˹W%~��^���#�����.w�:���"�e&�=rS!}���adc��G0��-&��W�w� � �$?ΰ������(��x���8ؖ�I2�*)�5�KH���x��|a�/*�����;��&�rJ'u�l�H���Tɳ�O%�}���߱=i�f�.N�>�xr�m��n
�26��>�]��P4�
I��n} F�kp{�5�e��"���� a@4X���4),.�/�������#��.����Y6=��<3B j�w������n�@0�2�'c����"�W.��!ve�4_%�d�!Tڐ1B|�kaU����o�8��i�RI~��X�BX����c�Lj�%0�Z��]�6��z����2���!�HU�+�1��f��0�)�#�B#��h� �@�=D> #߬ �AV>vr���eC3�з��-��#Ѧq戅�M
�Z3K3�jߛg_ !��	��kC����m�5�X�	�XJ�����*l�H1�1s4�xl��o��ʠ�Ɠ�0iZ���s2���챧S���.+���Hsʬ�s�:�G�7�b�pӽ;�ρ�Dîy���O�r/�,��m�]���Q5QF�0�F����I�2n�BRH���*�S����y�q}�Z��8ĩ(+�s���}�-\�B� �񼓞l�
�y�z=\�&��*%�1H�R�cn�Q5R)'���A�� Hk��jH!��[V��X�?��oYI���YI���yE6OH����*��T�O�ˬ��fӔ��9G��iL>+HfI�R�Y�1�&TYN�猒��,���P[�L�~�P˄L�3�#�q��h���0�#&I�~�/^�!��b�X�w?��hB2�!�Q7�Oh��
��1�����ӊ�AL:��]X]Я�r�W���v��m���̺�����bע:VM�j�9�]QA�	Wm��M��+���p�ƽf�fC�m���gQ�,�������_�Wl������L+s��M<�):hfO���3��4��ӂ<-X�6��EZ��9i�S�Y{��J�Y�|4%�*��L����y�� O
Ҵ M+��f��b�)�T��"�)��"�I�9�ٜ"K����d:%�s�,�u�,�)�\ah`]q]Q�Z;X��k�~�͋wp��pG�ywJ<OѩA�fVZ��9f�������ќ��rZ�z�Gi	S�8����C��4�ʵfe�Ej��0�س�G�����ze��
;�_�����!^������BP���eؒ�ZGW>[ǰ0���|���ᫀ�����}��x�Q6���ӈ35����OW:�e���7fYF]h��b���EE]hfYF^���0�2����4/8�MV�%YV�fI^�yQ[j�B�gYV��%�D���	��� c�3�Pۈ:��d��$�bN��)�:���	�R"����N�,�g�1	������Q��_���Op�O�+ؽ?c��k��3Y����~n�PF�V�$�1�o�3�;C��]�eI*g�n��+���G)k\D�<�RYX�O]�R��Ԫ��"�=�y�cV�StZS��Y�ÚyO�x�a��JB~<ʹ?4�1�~�+�z㋸����o��!��C�q�-@�B�9��ݽ����7��N��5ߦn���t�bt=~��nR� f�x�����v�͵���Wx�Z�� g��>����v�KP�lr>��ލ��9�f�k�c��
Y̙���(�6IgG�x/�@&��� ;ކb�����I/�s\D����s�]c�%��e\2<��s�cF�9R؈��>i��H�K�r�s^RQq|oL��c��^W����Tb"�ޙ��̩�
�I��3�D�2]Z�V0Ѳ@�%z)�P9+yawƙ��h$�l�oI���g��4�~�l�� Xb�#I�������7_ŷm=��[�{��ሺ6(�A��6B�j%�E��x����a��g[����.n���nb�wa�	L6����C�b���'��C~����7���?�3��;o��Oނ��t���f���ޜKSnt�cY5�y������]���d�{D�{�t��tZa�!��O�n���tWFh����Wb���%������r���$iM�T�iEm��U�8�U�K75Խ��R��d#
�l7��/��5 ,:؉��T;5����d�5��#k��
Du�T���Tݔ��X�kÄC���je��Hzǰ4DG��a�����*����W�r�����kV���-����2�̚e�hV!�ɥR��atÜqz�i�o��[�T����D�eq�h��-[���k��W��r�������or��#��D��);{C��������}>x0�O�|o�w�l��?f��dڦ�e��+�4i �M�QC�n�ʙ�1�w9��l^d�Q΃�������&�&$w$���!���x�ʸ���E�,���
�TT�%��9��)fj��qfi��`�v�P�*FC�Y�,I���ŞK:r(
CY��UE�j2���Tc��ǭΌJ|}l��č!L*�a\��l�>�Y�l�"9^��_�+�}Oy<���?|���!i�cI�D�U�,'��f�����<�0y"'���_��6�j�w����o���>�Ge&��  	IDAT��bh����\ȥD˸������DȰnI�l��t�c�H���lw���d��|<E�\B�et8�pwq�W@���9��.��Fݝ���b��k�������vk��q�3G�n\fy��i�f�w��a|<��.��-V/���Z�q@Y8 Z�!0�nWfԳ��F���>��C���ҵ��Tk~4���`���,uȃZ��7~����_������z���������N�ǒ�"4�	!�@Ƨ�wϲ^��A�H����~��������=��ѐw�~���!�˶O�U�h�uY��e�j$HX87��.�n�Fk�<q�ld�$H����n� �i3��X�� ��M��g7aPBH�V=b�I��
SW�z]��w���O���p<q륗X]]�`PJ5�����+��������~����];����X�MRi�R���H�������mS����7'�KY��/"_�Y̅u/߸�+7oP�������?z�c�Ɍ���@Q��Rr�fQ�*m��[{P͘׆��V���I����k��5��?�:��a�RI�s���2�&���Z�eNt��]�*M�6ϴ-^�XscLK��x�t�1���lqt�.M4�B�^K��0��@��|a�h�}�q0՚n�������o|�q��=n�z�3gV��'��G3�N�������K~�/�2I:o�[t}�`�Һ�
E%4������|�ۜ�k��6=�9������d�s�%~����~�Wo܀*���v��?�.����!o����9���%UK%�A�]��s���5��#���5V)�䜰1c �
�G���tN���<?�s\�*;����{�O��n���(׶�� �=��]�y��k+|�#��]�W8��C�NH�����w�=�~'��	:>A�{>���/�Qev���vl�mc{>R��FK�=m�t*��t\_�{��������:.����.���D��ƒ�δ& @Z�������l�I�h<e82��(�F�P��ǯ*����FjC���7OٓQ�BP&�9Z|�<�)3�l��(^z�*?��/E�V���dXʦ*[� $��Te�e7�Z��U��
K5@H]WTU�R���]W%���l�jeE�F�Zٍd�1��lhX��6=�n�)-�r-)��Y�G��|��O�{�M��#nߺ���*�R��|ν����������M^��(��Z�O�SC�n�.Zd������??��r�>���Z�7����3|��/r��/q��:y7ÇTj6<�O��6G���f^fT� ��<~���-�A�Ty3>H)��m9��B4,�0`0�b+��Ue�S�u	,�`��TUٌ�V#u�uM]7T"��e#-V�|��j��u]�D��}�^v�Rv�i��F��vM���o�_����sm|��h���ׯ����h��|>g�F�c,�����Y>{�@���l�	"��s(EE����Y�/�'�xK
�y�$�u,>>��ޅ�̺�1EC�$�4I�p4�4 ��M3pz���g�B��G���]��N�-:
}�n(9�7�5�������_���2��#�З�_�L0�R�?S��_Gz=���l��X�s��h�W˄��r�u�*�xr�5o�1�y�_{��~��cq%�:R�ё] ��������"��mx�\l��V�o54Y�ϐeEK�ٔ	�p�/h����=�m�V0�y�E���->?��'��)k>;��kK|�D�������V-v���}��q���O�MGh͡�����]|eវ����V*eq�l[�>�e5�P�2�'� b���K��#4��eR��kt�[t�'-�<��'z�S�{����ˋ��������O�ͧ�7->��l��FH)�q�����o��zm������c@ȧ](-�r��+��R6����iٌ͝�u;|k�2GUH�+�S�'��S�F��&���'N������I*�	��F�47߸6���9�:�i�:O�O+��I����M���>�7�/�j-�tcE��1����������3��u�18�"�
d,��v)�jY�H���X����-V��J�qڰ^/*��I��f�P�S�Ŵ�CA�t�'+�c�{N�	 ���ȕF�a�hx��ś��&��F΢�x��_0B<sN�&���v������R5�9-��86��"�h����_���nT+{"��u�Ƒ9�Z�y5��-��4�A,�]��|��>�u�?]��h`�q�k�;�MbtK��0�-@���6��!e�<��ihLO����>h<ЄAk    IEND�B`�PK   ꩈWQ�O�  N�  /   images/5c74bc75-11cc-4f27-b1b5-62f572483d6f.png O@���PNG

   IHDR   �   �   +��3   sRGB ���   gAMA  ���a   	pHYs  �  ��o�d  ��IDATx^��y�l�U�~WD�s:���pK���P�@2B�F$�~~~�i~n�׶���1؟n��ã?�<��M���fh���)$!	�4R%�J5���{���{G��?"v�<y��{�U�w?�f��ܱcG�X�b�Z+DU� �{�1��"���?��������+#�]Z2�%m����"�W(6k�?u�B���0���_`�V{�:��J���И�GsPeXT��=��/Cӕ��� ���S+������w`"��)<u�j���H�����g���Q��E�E�D�H��4Y��C�*'-/G�K/;�7���Nk�TS{���� �^���B1���@������w��O�(���"�J�������� ���Ù]a��縲[��R[��P�{&]�Q��`T�ݧ��k�\hLE����;l=�Ȑ"
���2�;D��Ld����NéC+���t��n �TX�s;L�GIO��N��"�D'lO�������'��1P��2�o�u�CADu����>���n7:����y�9�s�BQD�V�M�?������hȰ��Q���(�U����e�����ɔ�����z%R�a�,EYmE�*zTP:l���R�)J�445P`��5W��B��ad���s�Q�^��K��gK(�-��$�>ΖeEQT�e��_�
lI��x����b4D���ɲI,�_PY����� [�u�|[.P���P�qz��;��9�fs�L�2���saX(J\>9m`�Z|;Ň<&(����-�!���!jC�e}XR���mQ5J�b����1�#����a/5��)Z����a��i�C�G�JZ
��QSRc���k�zS,+���A1x�������S��\;�4�&�Mj?i�j�J@�7�fBO[z0x����dyV��J�'�#ja�$��Ĝח����3�D�j���*37�$Me" "I�/��JD�A��˓E���(��JL��)�J7�4F���b����d��Ո��iS�"F��'J�H4�h�����fӫ��i�Fzj'�`1�`0AP,bPcPQ�D����FP���T=�����58�n��	�v],I�qA�3�g��kn/(s.C��OH�x%��:��>Q)$F?�p���kҥ�i�. ą��b��HZ6�I#��=�￯�}�!G0����c�nP~CB$��<!f
�$�#F�_���2"J��1�1�����>W�1`�H~��K����!>�x~��A��*��fْ��L6�ĬL,3|<�CDE����|i��,�-�1�^�DUZ�_��d�N�i
4�0�t��1�N�����&p$�ŶѤӒ��̙��"��i���-�/>��4iڌ*I斩D4F�ƴ�i#�H�>$ɓtռR�#EqD���:C��3�r���S!ҧ��靁�����5Q2���A���Q�Ac7���P2cE��ŏ�C��iQm>6E��~�S��9�C�^��dD J��H}u���h��Jz���*�.����u�cՖ|�U0��A��	�ɪ�F�X{�sW�4bb���!j0! �8u���:$&Db���D��^���c<6l4����F�Ff$͕+,��� ���"ZT�.��F	�"o@���=��cx�>?�Ib�c�!k�"�6z�≃���p�s>�r���b�˥f�g�=�Ի����&�=��W�v���T��ӧ��'��%Z6C��ز��6L�c;I�#vԕ/iJw�W�'4>p��k��	��f�7l��>����m b���l����ku�d�ύ/���z����N�3����o���Kv�kT�i�s!MkJ��fR�\��	h4@��6I�*&n��Na�Ê�%���&[^۰�W�r�ק!�H���٪2�h F�A��'�*Ƙ\nHbR��aѶ��(&��O+�9U�W�7S���g-&뮰�Sz
j���Z
M���/�{�1_��~i�Ԧe�V�ŏ���9%M�M=ee4d2mp��ش����$����m�	�|PL�C~����*N�^�O��`j�0cN9�P�܉���=���	i:���M�s5��*��9��4�r�
c��6D#Xg@/1�Ⱥ����͜ג����p!�P�HU�h�g��ՖZ��Ֆ)-�oh��z���"i��yI�.�Z!ZAE	�~��]�L�(6i'ňI��˵1�N�~}T�|��l2a7N��|=%����uʹ��>*�I��Q\P��K�fA�����}bi_�j�vbȻ1���%�@kӶf4�	�E��#D'����Fr7+t��5K�(�t�N2�}�_Z�EIk��ؕ;_��tE�� Y�N��4�3Dj�>y&�tGR�"����MΙ�7��̩�C�[A��F%=]�f�3ߙn+�����T�i~U��*1�7�Stg~�ʙ���v�N!3g��+�#9&͆8���q($�8�<��V�
P(Bn������BǭϜ�1i���Yf��N�XI"r�k��&7�<uB.�݊ZI�1Ygҁ���V��~�M���g6�|O�1|He���Kf:�T~W�dc�!�ac������}�8�(�s��5��2;��w`✴�V�Ě'�{_��UI��$X�,򵚙h�}z�1f�CicZX9M��"�<U/�@c��<�4�i�BaP��^��GT�_ص;&��C�������lv�,��i���S��	������v_:w�p��$����B,��PR�B>�}��R~3�6_���q���M����/,�ᭇ�}�I�E�(�
:��g_G:��RQ�P7Ew�ܪRxp��AgR�N�rP�<�8�p��^lbF���N'���3�Kg���ExQ�_��$u]L:�6.ǭϜK1��q�d�V����	lr�E�#���M��4�h��Q�^Y%��Nw�t�����(1�u�&�9����B�Bc�9}���V�����%����U�D(����4�_#���8Xn|q0�Ja
V���)G���L2IEO,"Ct�=�U�D��b�R��P;�J-�"���$���|#"B�� ^p���Ka�)(]Aa}SQْ�)�wDI��(ꀛF�I榴�I-�{�[��Qͫ�^+�7e:m(JG��?<O�EȦC��L̨�1����w�[�9�B!(l�N&�]�d�Z9��-�*�[�{vfI��N�Iۈ����0m�^�m�!�r�	[�QY;{��mK�ION�$�AR��uwj�"[%��}�0g��+0v[�/����`u?�4�Kӛ���1����uܙu�~�I�fy��ik�0&�b��.�G��VqAQ�����}����O�^r{b����3o��z��Lj���D�U&�cL48kvt��WX-���;_�*6��ݢ�O+�����^�I�����ˇ�-͏�W�6R����P��J��F�A)Q�+�G��i���Ĉu�̙YdV��P��~f� 倪I1�e�)&c�>)U0�� "�|�"����@0I͠���)#uJCi�g�g�'�7�a����M�ՙ��SQ<��;���8sv��; y�$R��"=1X=5I
�5����)��`$}�?�to�ˆ<�(pT
����,#A�=�L�A�l�mj�����dHN��3���J�2���&l�s7 1o�.�8nq�<��m�9��-��]��V@b�$]s=Ę�&/�$.��,sl~��d�}���e�B�5��f���箣ӓ�	�[_�̹�#�LK�]p��?�	t�μN��͖���E%�_D������ɜ3h��"�P,R���)�!���v�B(@1���ndڵ`@�t��2n�(P ��������H�3K��J�n�o.���]�������R�y�e@�]Z��ߩ5�#S�ݚ�bz��i�r��Lb�$[�nґ/A"��hJRv> l�y�E�Ol��f�E}� Yj�P|^����K&��Z_p�"`��]f�5휋���	�E����D�hSl�5�C��해�"��AT M�3�T��e'�ӿ���%ݰ����AU�/'
U���=u���\v��fN��1�_��ZL4QCkJ��MJT&:�qlG�U �ĸ��2ŶkT44���!z��xZ"��cz`+�8�1Xk��`�a�����!W5K�Jld0ɏӃ�u�5sY�c���Af�%}�>na�\@�KCJ$,V=V��Px��iO�*��`�GD0>$�,��<���s$`�К��{�hs���jm��}�Ӿ�S��
0H�5�%I�f�͢�"1��,��o�������+4�WE$L$�Hhb��6�!��vJ�L�0�m<�����sYː������0e��z��c_���A
S�����$JJ�c\��>Ԩ�¤%Ė&Lf�Ŧ!���|Ӱ�L�G񳔭��V���[ϒ���m�C�[W ��Y,v�^�$��z�E|ζ��_�(<e���Tw���.h��4ʞI
���KW�p9�r�
up�0�-������� U_M^�Ŋ�{�W�I&�g���%��K���aǵ��-+���I����!tq�G�k��~��I��s>�͇��_t�/�$W$Ő�J�5i�K���$ER�9 %m���H�E����&����3Eڮ�s��;7Gڪ��Q��[�*��3�E�ĦhP#"!H9�:�4}qL떦�ַ86�:� ,�8sU훂������F#��D[vc�$4셆-�ى5{~�n�3M���аZl�Hv
�]z���t�1P���0e;�LC�4�{��!k��>�f,[����}�*u�LB�n����8e7L�5�0eMb�^��iٽ�әM�l��ʜ�3���y� (��Հє���'!���"LXQ
"��I��tC���ϯ�I"u�"����n�bM�JJ�}�4"��yEz���Kh�&�Sh*ߩP�bD)TqQ)b�FA%J��\�u���V���Y]ٟ��хѦ��Y�Z�^�n
����.���)b�ӄ�4�O�&��BJ��IIԤ�nzM��(9_t��C��n҅g΅ib(�/�B�;��N:���!J����D4���hj�5ɱ��\B��sӧ�?��w}W�ף�]�4MC�G|��l?Ѽ��a��[��<Oi+h�MO�3�L .z&��J:�2ʁ���䙟��u����"�d�� Њ���|�(h��J�i*7�\�i5{��۠7�.��<��w�w�CB�s?�s|���m����H�*R^�i����W��k����[�ŔU�@Xµ���ׯ�P���=:���"1�n���ƕ����z YM�\|��z��;�P��J����\�=��/���ۢtiD�ĴP\��˦�H�Q�~�������ɓ�:%�EL�7�%�N5��Y�u��������e�^���S���s����uZ� n��/Wb>�c�Ŝ�5�/s�f�+�|��'�ʟ�%�|S8blQ��.)�"T0�P�WWW1���n��6F��1i���a:�m}���ò�j5�*��Y�dw�������O��X�Qt#��|��;��0Kʛ��#��X,�F�͵��e�+���}z�����A��GC����B�?9t�Q ��:��T҈ v&㮳;z>��Vϸ�뎃�x��Z�\���/PB�1��h���HReQ^��|����\���O?S�>/W�P�Jȴ�R�E�B%���A��u�������5���B����Yf�%�1O����,rU���\���=O8bj�T�2�t������7J]���y`�t��/n7ɜ�K�V��(Mi/\�B����0�$��ZT!TQ(U�0��wJf�L@��j�4�l!F��	�R��B_a��RX�Py�i��$�&���8|�|QMQ�(��0���J�g�QTpy%�JR�@�۠�� �Q(�P-�RC�^�G��T�E�(1VH�B�����U(� �6��2{E����c���.A�i� ��<D�mNX�*��gPG�u�?��T�#�i�?�Ǒ�8R��Ɓ)�I�@LZ���#�c�\�N��DX�s�O-�c�8�����q�v�V;NN���k�(6%�2d��A���C�-�{�f����XVk˪����i����co{7V��jI{*P�+H��Ɓ�X)�-�*wNN�+c֫��ö4uˬ�h�ɯ*+��F������DX��DS2��r����~��wm���U�����������d��$*�&��D�Η��?�/�rv�b�Z�8�t�w�V��w�BO�h��>+�Ybg{_a����f��M>�<yz����9l����;(W�Pg�JW����(�+z�*�+0�ɠ:�.X�m_v'��u����BzF��|�Bܙ�<�,��<#���e0p�
�\g���u]��iq�~h��9��0iӱ�G�G�C��C���;��l�˿�K�>��T=��p؅�E1��5�{s�S�i��QM[wj#g-+E�!�j���j����ui�(��r@�0��tJh[l�"�L.{(��nJ3`�:�K�qTT�M���Te��g��+z�&�o��h�̞���۫VJ�H,��+i��Vs��~L��!c&��
ezb�X0��-��!+R1���R�vǝ��DU����.(1�vPe4Bo������c�����
FްZ[PK٦gH�m����{Ln�cC����`�*�e)C��:T�i߸�J��)�`��rgQ�B�M	X�O5��_��O���>��>�!âb�y�[��y�:��yE-?ZP�t�A���8/��2KK���'��M�$I����n 
�$giZ�Q�EC?
EPʐ�����^ݾJ[O�a�]q���)��(�4��p�^UPb��T��Q(T��*4���0��`΃0&b����>�T���=K��u�)�8) ����p�v�a����N[��VO�Ҩ��a*0M�Aڂ�y�U�����Y���7�b���`��v3F��4i��1L�6�I4�v���k��M!!1��U�ɍ�g-U�h��MɤpL���[��n)�u.K%C�f5�G�)mz���W�Ah���u�Ǥ�+�]�
&;�v�G��]tCx����2�$�Y��J�G�K��)�k�AU	���\k4
ycR�8�hQ�+qrڈY'��0�K��'QP�(�Mw2���6&�/��z�yz���$�gz��}f5B;K+)�H�t�l�HbR��e������T�s�g�n��
��*BO-N��9.���Ǭ����@L��y3� ����e�ύ���v2a�-ؔ���	�9�t�h	��`���]^�*�o�ck�@]n]j`��6���H��)d�K�S]�k|�F9�;v�4�õZT�j�]m��6)q&��4_�YH����_�Q1A1&6���5)����l����1�|p�6�.$+�YN�~�t#�z�C�� �7��'K��:i�u\6z�]9s���G:���Η2�v$4/P�F�����s����~]��7�<LF���ZC ��>�X�3�DP��<��� ����.h�b��V��t�:8�0���h�)y�(3}$麦;h��~n�9%��?��F8��r[�BG��͜2��f�1�K�zdNbJN7���>�
{��Z���.�ؐ*n�X������LI��ZR��0G��7�ԙ��[��q���%8=Tv����6�� i[��	��ta���fS�d궒�I�HAPC��-Y��G�㸸i��9�ɘ%��Ջ~�ס�I�<�f]4���J�ޏ�/4K@����&O�m��a_W�ь�������ʽ���I���������`T����!t�
�W���3Œ�!}�W�g��^�5��:�yQ9J��2p�>��'k)0�ٲ��T/�͜���&�!1�-.*1����\�iQs#�s���ڨ�M{��Se?������&&Y���=֋6m�:���$(-$Ǖ��!���ђ.Ef�*��h��1�)��&;���D���w�!e��/��H��EA��lp��ǰ�b�}�b�]��'r]�"#*�,�DACL&���1z����95��������S�H!%a⩧S�-F�v���CS�S�r�Ŋ��#J�`�l����IQԘ��N�.W4=Q���HThۀ���B�� uDjOϕ� �-�ؼ{~�%�h�<8�#�'�0!�odK�����y�&�����aWR�M��+8c6�������$�eb-�B�`Y7�f_*Cj1�h�Z[�mKlh[O�v�GS�zB�m`:i�6�Ht��S'X?�"�ڳ;�C��Z&��(w�k�X��ADhچ�`DaK�.o��x��^�[��V��ַ���S'��t�=&m���&�fgZ�5��jkv}��z
!`��*���1��ȁY���H+�sBS�LCÞ�40����h�����u�tŐ쎖4+�e	�*�	>��1�U�V�Z�U��G��'U|�`��!��.�=�c���M�=��R[Mք��<P;a�O�t4gs~�}�-�TLB`=X˴�4eR����r]
F%�F�K��9�>����ț��f���c��5_���W�n�Ř���<nho�m[�^���U}|�q��{Y���+#������[W޿~�6����z����!��i��щuڵ�:zJ19�-�x�t�'B�k�K[8�F|��9oL�}M7r>��
M��O)V�$g�g	GA�F��)W���j5�e�r}3C�C��3��:*S-�4=��Uli.���&�a������I&�X������$��$�dM�r��-�\L�.d}4U���?�q0���=�+��co��n���O�~���/���1&Y���~l�!`���k�>o�#_�KjԧA����%�lp�̋x��|�º�7��&��%%��15�^L� J��xS��37��ԭgTU�ڣ1`�"��oJ���C!��zJ]\a�� rer멁I���c�
�-MӀ&y!Wd	;ϟ�I�E���6sF���%�K�
��1D��/*��d	2���;x�rT�����fZS�hR��n�D�tR�V��gIf�K\]���FA�xx�����x���Dxы�6{�=�.o��G>��?�a�WW0�bb��n��͜�{��)gϞ�k^�z��E���ԓO�3��կy�z��������O���_g�m�XȌ��vH��A��e'�$
��ÄH:^���"L2�d0Y�4]�(x�]�X�N�H:!ͦ�n��g�
�@�t��ɧ/;U��j�kӢ:�0^�L�{!�8$w��H��駦[���#�)D���d�,��FV��(��������ל����0��_�Z�}/���K[x�|�C�}�{/Uo@eKbȺ�8s�*��ӧO󶷽��︃�x�O����������Y�����5�y���esFaN]��,u|�4Q�`��_-Dvj7�;����Hw�����d�N!��H����젺r�t6_�ԍ�i���w�r9�K;$����1P~>�;�J�y-��9���=c��˾&D0!툌W����~1�.,�m�}���'����g�w߽�~�휿p��C|���:Ǡ�/Y~��p-A�4�����׿��ﾛ���ԧ����n��[��ӷ��W�Į�E@<h�pLҀh�,�H�z�P��i�����QLW�Bن���N���ڧ�!�ENݿV��P��1�L^��M�n�"�Ic�&J$��&��O`[v�,�$p�+� I.o"��n���Bw�����5_�����1v�vy���8y�$��ʯ�%�ߏ���9�d�#>�`������x�9��s������uo|#U�sSP8��������7���YB'���׻� �}�t��t�ق{�å���z��f��V��r�>u�=��"��4�*����'OYTc8{����_�D#���N|���>s;��$�q�l͵�3��p8�(
VWWy���NUU<���|�7}ox�ҳ�d"�\A�e�#Z���e6���0́���&�w�uX��-Lzݽ�1)��^���a%��E�?�M���8ؿ1*E�(�r����~���;��gϝ���6��w?����Y��t:]�rd+Yk9�<u]��p��	�|�I���7�U����Wy=,$º&ͮ�{?�N`�8n�eX���qӕOXl�E����� ���k`>�ϝw�ɷ�����XÝw���m�QUVWW����%�b�'O����&����6��~;'N�8�9g�&cּ/ֵI��ߠ���b�����kB�f���i��<�]������M/j��'e�mGf�����S�}�Yvvv��;9q�����m�tj?�9�1loos�wp�w0�L����
^�W�i�K��vS;,~{,>�ɰ���t�����?n&������-~j���3]o��[����8W����7�|�\%=O�v�,�c:U~����kC{���CQN�>�k_�:67�P�+++�eI]׳��.Q�b�#EQ���B۶\�|���Ξ=��^&�dc���蒏�b&%���ܕ���c�c���5��+5����(ݘ��Nȶ����F{$--�Z\t8���7-�N�u�0�����h��Y��%Si���D�QDRQwU�R���j"j�`"~�ui���^���-(�� 2[B8���`�eee�~�@Q8�fd��R�!��!�9���9{)r��N�k�K��(�k�TSj���d���<|�9X�Ds/u�-�$I��]FR�h����cgF���Q�dR1ٙ��d9�h����͟j7������~*��;��$活������iS=T*��a*w��צ����?�|O,>eg�RUaƈda�I��JN�G2�O�҂��`Kz��g�#��g=ITڂ�T��������RX��>Y���PR%����L*��9��ye-C,���bC��is���ݸg��TRठ�E:x�V�RQ��R��7��vbb�2�"[3�b��kSى���)(M*���:�149��������6�Ai
*[�r�VǤgR�`,+yw��k~�#��b�Te5��u+x����R�5ox�����Ο?�<��}뷡$�i1i�)���O	��o>��-`p�%&��X�ޔt�O4�)�W���:�Xj1I2@QG��.�D(,�ϊE�s�)N�)���E2�wߩv	���7�	;l43g�?��&��B"m���!qP�!]�Ѥr"����Wƨ�D#�A�Y�z`T"!FBa0'W��j��^�mҘO�;Sd:��IR^GF�$?}�v/�oz_^���B�s����?̿�����；'�x�����e{{;���y�s}�|��y�;���+Ws~۷�-BM��F��xF�G���G�`�v
m�)�Ҫ�M��B�۵Bkm�P�<xz�*�mC5k̃�Y T[��,4-e�o�C���q�;^�
{�e�%w�#Gm;�˜�wVOh-TѠ�0~�6��Y��lẋI����vB�ewc�X�9Ch۬_wea���n��g`�갢T�n!�D�8�Ҭ�x�KiK��ۤ�����ĤCq\y�9¹MF5��T��"�4mK�/A���w��W�d&<�S��?�����Y��A>��O��Cq��U�*�i�9wt�T�^�7�u����\�|�D�"\�F�
\���I=��1t#��b�U��g{��[�n+({8�ģ��UU"EɰWѷ%'\�ȕ�ؒ^U�Z����~QR�Ʀ�0=����>,�q�Pڒ�-X�R]{UŰ�1�J�e���1tF�O�b��)@���>$3���Y�%U1�?��!��b�z]�aU0�J�Uɨ�S���1D��twS;y�(���
�X-+zeE���W�{7B=���~�G��@\l�y	�0�N��ކ����m��9�?]=?�ɜ����i���8y�$O?�4�<���L#"��܁��c��#���KiL�RZ#D�Rp��-��X5iz��H��)��|��.��%9>)���ϦT�A�%N2 5�b�=�JK:��X����xA�!ZC�]����_;��hi�b4y�"5���$�CVOR4��xB^�@z�n�QR3�MZ@%�%�Z,��(��&�1%����۟�v�/_�G��3g�POk._�L]׬��/vG2'd�=�٧��d_�'�|��W��qe�[�6F��I�jҚ�[O.RHF#1�a��������i;[����T�7��n?8��+x�g*�̑�H!$��Z&Fm��%��"!�<ؔZb���hMns��vv���*1*]�� I��k��A4B��:F�"�5@^yCr��|j*�}3$�I�IL�V�����(F$�c��D�!��3c���Rite�
�z�Q����s�غ�E۶L&��e����1���B��?�0;;;�v�m|���hM������FM�p�#�>%��`�b�A�f�A��sC,�
��j`I�I�3y�e�/BbP=$%�I�N����"A��E�M�D�3�B�Cp�U���Bv�KE�wdZ�H
��LUF��$�EfzG�]��ڜ����y= �_�f�Zz��x��l�%馝}6J�I�J�����������2�(������ˬ��1g�}7�_�9�4M������'��~�7��G~4;}t}@�h�@G:0���&��*�Z��?+n�9w�v�2��9����d	̘M͙\H1���,�f�tx
051y��"HI�<�B�`?<����NO,�OK>ZF��5�@WAQ._��;�l_�f��)�~�Y�z�I��e<�4����5��{?[==��|���e4����?���?�QL����J�	Kd��d�+�1~��Rk&VJ��p+/�.�13�}��bF9S�\����&e�%a��]]ٟS,>�t���uC�fn���=���O|����/~1�{>�اx�󬬌���L&�}���d�UUa��ܹs����nj�WV���_��?硇�&�z��1���Nǡ��r��%XYׇ�����s�I�]G�n�# yO�����aмW�)=H׎ik��'�󬲼}����q�r��?Lm���s$MQ�<��~�I���x��y���1�ɏ�O=���iM�4�z��n��?Y�jғz�O<������.����������������/�~7�1 ��k�������}�:I�R������э�{=,��8��|�f��94�S�|�9���uytQB^�fϕ^M������ӟ�)��?�)��9{������{�C�B�NU�>.�u��%���'�z�w�ֻ���dcc�����]�����O�C���gy��,ӵ��},J��b�IG�e��"���2�S7������&��EN]�̦��p��]�ty�F�;є���0;�u�w��|�T��Oɚ��_����:�R=$�F����3������?�Ϩz%�X�y�=��p�w�λy�ｗQ@QU4r���b�n;i41y������+�އ���mFkl��sj4�ĝ��?�|��L">� y���1�ie�-�#eע3t�d~��Oo$2͡��(�(�MK�.�_+)�z��F]摜�w�c$4*�Is�W�Z�"H�C�ڼ�g%����%�l.&ͳ�SG������4��".[I�>���]Y�t���2$?N>*EpQ����5��O���c��� �g�lp�*8��{�YY_��G>���W����}h�lno3�L�9��.���~��~��|'�<�EQ,��d��;G�����>�,��^�O�p���t8�9����0s}�>i�\r<s��"޷�>��O��AUR�l%�Őm�v≻��Ul�h���AN���YIa[�$�VW��� .?�ON����Nvas3������3��UO��6���4��ud���5��i&�(KuH���V��F}���tn��L�����{��e�`��A|���Ix��Q��)�U���뗌�)mlr�[Z�V�u)��$LSb5ka�Y^%{��1�[;��p�|�<��1�kF�>�(�UΙ4Cu�Vn�#���y���Ac�hiڦS2�}/Wn���o��8�*.�
#�bQׅӴ��gl�h#+����Q��'͹)S���4��L�jl� d���}��N�(�,h�lY�%����0j���K��!6gjSR��n�p��:F̩�_�?������t췋״L��0M$�@���3���y�#I{u���L��b������.�����{{���2�,!jNKg��{��?�?���Oqi�2�z�+��aU�*��"I�c��q��	ia����!J�<<퐯����|O���ƭgh�K#��F#P����@�3pN���S)���C
<����Ġ*�Rzg��AC�v��K͠�x����xw�+��S�y�8cB P�c@C6�����l!:sǷX
c��l����O}�8O���x�H嘄6%?���O��8cSB41�(�AL�b�3'Asm�61 �����e>�C�W>�)�?����oXY]c��U
W�\��=.sK�\͋���P��!��T%bS?e�7L5�xv�s��	-8K��/Y!ώ�3�$f�i[����ơa����l��mي-Wۆ�ز�l��I�i�gZ7��g�e���5S���o�	-{��j�ٞ��a�8��~'-��J�$�����=&���o�Ě��e�g��	-c�c@�{����4U滤�ٹ�S�D�-<W��r���l�)�~̶�\��l�S.�)��t�4ǱG���`o:�Gp��I�A�:�a�TU�ujV"�168�����I��Uz)z1 @�@�P���;���
�*���RHJ��$�L�pkR�¤������9U�A�_&��Th��m�$����\4v	!19�.	�c(���PC�C��R����=�D�� ��Dv&$�����$���쿏b�t0&%��rn"����TXŉ� I�@l���F�5����Yj��>|7��=q̬e��L�I##M��lg�d�t6yLeH��%M�>�9`Z$��*'?`Z/V���M������	�%�b�4���|����`�����~AG�ߡ�:�4]`er^6�������-�ȇ%85�JJ��#�����LAY�J��"�"�^�����6��¹��t!�G5�5pS̙�nl޷<�܈s�r\�����i����V��o�1�������㐲 Ki��.�"�N�'�Oݐ����$�B�5�i���\��c.�󥘅�h�*0ɫ�,���S5��,EH۞�J��D�%��s�틬����4kːO���sB�*J�)�{)i���M_�j16����܊J$F���$��k�Fb�%��%�	s_-r���!O�$S�Z�v)}�XMC!3����@!��3�m�dk׾��c�� �n`̪��*�Ȩ"&�J�����)��q������� ���mf�n}��3�yg4_�1��fE�.����ق���Ug�o7Ŝ�[���&G%&�(BZog�URǆt;��8]�Bn�#a��@��oQL�u��iv�.��Z��I������Nr�3c���&��Q�G�t�ɡ4��As��ZshQ�(��T�6�,�����Ƀ�td(����8dc�Q�ȍƀB�qD��kv�qpS�������/%�/~w,����L8�etL~�-���s�)��t��桒�q�"K����6�(�����3㐅B3:�V����6Xo��YI��/�wyu:o'ݻ2�t3y�ΙHA����|��ڗ��K:���b?��+H�u��@�*��!uP��k��^%m[ڠ�&	�h�F�"$�V�5�S>$*�k>O2����M�{Ǵ,\܎KM��@��3&�>/ހ��%��9���m�7�T�4�.��]p��{��ȫ�7͜�д��C�|[�*�R�HiqR��kJ�-q�ĸ*�lY�ڂ�t*���e$�y���Pz`����l�qF
������+P;G�8����;(@ ħs���bK��pRT���Va/
��TS���$rY�K�1��4T/�9<��7�??u�p��(楦����I�Z�M���g����Z&�/[���
C<`X�8Sbcĵ$ۤ����6���\T�--��Kq)P�;�~��;w�"ť���ww�`���[^x�d��d�ݙ�wl�ߘ�����;�*p����b�DǞ��s1��=>��0N��47�⌊(U�&�� '|��6�L��_��0�(����H�@0�/s4Mu��Z�.���Ĥ���z��̧�g9��n�ɍ��'X�'������)��ۓ9��^ +�W�H�X^c��:���@&�FoY�����I|�*���V�r*�c����g��  �O�w���s�W�$Q`m@�d@wT�P��LY'uVgYdPų� *�w��\j.�n�i%��Js��i�k	��2Tk\�=T��%߄b2w��QO;���ߓ�D�Z9�8�g:ކ]�x �����B�C��B*�!����*��(`��6�,/XYU��iz|y}q��7��A�I�_\8%1�CwH�V٣[|���w�)�2�}۔� �Mb�4�]^/\�3%�)�����5p��Dl���؜s7qfҥ�:�gk/��{�Q���A�FЁ\!��m�+f�����@CM3{`)��M�^��V�r�<�k���ݎ����8�w ��n���)U����f��2�4$�K݅�`W��~-�19R���R�F�/k|IිCyd�
c��Ũ|��_,����φ���[��U�(��Y�J>TQ�:#5��3��VV��nMJ�T�?��=Z+��'{��bۆ�RV�yl/�K���9r�<9���}��X��7��"1E�����&_9��|=&,��@<0"X�%0wə<��M����`�sx��Mz�NQ&����ct\&�kK�p�A�ET�����$���+S�8�AJFٟcd8[���wn� ���o���c;8�Z���Ӡu�q�M���
M;��˗����"��6������n�>����������D(�;�G�t&
�MS�8Jy�~%�1���^��ސ�T�+����lj[e�m8���6m<��q���Η	�8G\�6�Z�cg��r�M�hS�0��@��ݻ�p����0W�߳h��y�_{�R< �å��}1׶����.Mzt����w.8��4�����ѝD�x�z4gV��@e�
eh{Z~��;�r��'���y�f�رO԰*!pbq`q�4�f��;%dRF����ds~L��x냟>m�5�)��]�ͳ�|��32�>�W2r5�Toe~�W[�7�0B'+*���JVP[��V�|C�o����
�%:�%��b�*�NJ�c�|�:������"����S���)<��s��&~MR֓�/��t즿�{�����M��ų�Q��IZ|uuI���S�گ�n���s����3(%+ڀ[�	�n���ҷx����J*�O�TA��[v�|2�a��(��Fxg��.ע+���j`����Qˏuh���hDR�W(�jɍ�9�M���_V�"�y<PҌ�B5D���F�L\�O��?#`9*I??H�1wJj/�DC��+]��5J�H(�4�r�+j�;J[? �r`V��Z<������J|B�4,�X�< B�i�cu���HND��f�e!��.%8�2�5Z��,���M�U$ԟ�QǦH���6��:�bB�8r5��N�ٌo�uN��h,������|G��I�-��jol�]�T�j�P����a*���������?���,��E�� �����)β���������r�W�w�m?����S��c4��P2�I����T?���:�g��e~��%�:#6!B!���<|f����ӵ�%E����V�_�8������|^M�<�_
pκ%{�x�c��&�֐�����V���d�խ�\+���L�p��T�m+ֱC���s��1��⒕Ƨ��
�de#�i��4_�U��7�/��to��o�
�:�^Nd0�<.�T��=Pf/����7��N���Bun��jHϕ������"�X�Y�1���+��S���	�!%>:~�ЎN�S���t�<ů�̈́��	�b4�s�C��'��s��R�/hdV����s����ӆM���('Z����}[��sאG �XN�%����y�q�bQ�%���8V�C-��	�v7��#2	s�mD��e,��,����ņ��~�o��)�\��g.2���R A��6:j���W�4���~� �n#���_Xs&��V�2����-��R2�_�Wp�L�MLc[�7v��8:�S�#T�e���W	9��0�Ir�V����9�b�}��	�����L�)\�w�d��L�)J@1*j0dN?�-&;lU��}ۅ?�zz��DNH
�4�'�bR��e08H���!���.<W�L�9o���!�p��9��=�����	)��G�*��K��^�	R6`?���z'���;(<�m:i?��f���F��|�	���3�����hC�I�M�lI,�uK�?gNeG�`��: ��=��?���p1	.��
6�����T���'�a�8s���Y� �-�y��͘�I��MЄ����u�{t��M�X�j;՗�Q��"si/N�Y�2	���
R{h���9#��j�J����������>�sM,����%sE?���N���qD8���]��#=jVy��fn�@��y�:��t�O��ȎH y6�/+)	3)vG��>:x���P����\z�_y�<J2�Ի&e�K�n�F��|-��'�S�����U#5�1YP&V{�sָK�O'_�	풞ƻ�-{lRuܟ�W�}��.�1�9+���ԣ��X,z�r�Ȱ|���cϣ��bf�����m͎+��2�j��럿MwyXqČ��� �fM��Q.b�9�E�_5�|=	�U&B��E�lX�X�����r2H����3���)K �[B�PQ:y��)�w�?[��{�6f{}�˯����f�4S���&�~m'_�M`7�)-�fD(��Ie碟|u��+�.�#�ļ�X[��T:���?��lr���\Tf󷃸HB�)y7]��E{����e��ū���ճ_�|�����Gw��Z�)��Y$Ŕ�-Z���_#�����F�%�]r�B��i.4�;��u�6m���f�����ۨ�ʢ����@W����~��Yt����Xu�v��v�0ۖ��z��i��'0G��␰O���\�4�d����8oMq��ajs�\��qnKצr͈�TuI��!2��j���Wb-��o'��-^zcs���!����(
p�5�����OH3"s��\�Ƥ*���O������u!}��"��{JHd�CQ��z-B������S��D}L�f#F,���Ȼ�np�*�*�f-��O3�/n�6�p9��[�X��[F��E`/WMoow�1���?	��\g����1�����w3�IGI#��a�-.���d)?�-=��1^h�5=f����X����Dg�q���r,vSU�Ɓ��ѱ�G��s�5���d}��x6����ӬU�L���FK)�8����lp���Ks'<.��X�%5i��K�ʹ�k���Z��s8U#�ZAV�.�l_�Q��q����Ɣr����yR[�[���E�/�:�΁Y�rr(0ֲx�x��$ Ll�(T�xB4�s�x�b�<���']΁S��²�R�3�_��u�%X>�dv8�e:�&-�zl�{P~6�����V�^�$4+zh���g�4Q>G%~*�Ϝ���E�Ϲ�#�
��s���l�Y�j_)�Y�4jeF��)���e��ѾH����R��7~PD��!zu��*Zu?�81�! �=��Q�Wܟe*���F�[|l8	�%㤲n��1@��pt~����Z@�f`�6�\%�ώ�����y��Z�Nn$�z9�_�PZf�F=5�j6�|�rQ~('c��8��%g���|�?�ݍZ��OOƛ`)�lD�c-������^ŉF++�#�sk<�H���_�9�w��sÿ>��~�Ntx=�������|�3�_������t���)�뢐@5"�hb�Xh��R+�u`3�e�z�9�۬�f���c�$@�>R-:�)> "Oju��x�1���2NO2���P�%u$$�P����GF"~��8�&�9�`��M��Vm�����\<"󵌛�P$u�:�8�T���z�ę%�Y�R�"��X��y-U8�#9A��?��B�������*��c/�KZr�/�7���G/�y��'�/�q�L�1�qQ��Է��Y��D׏[��*��.����ih1��El�x׿e�:�+[7���l(��w�)��Y.�.q�C��PSΖ�U�1�����R�\T��z%/9�Obs ��/ބ��W�SL�Y�Mfhyc�����Z֡-���Z��(��[TDi�v�k�%��Hxr,\3T^R30))����bSn�]��T\�qFG�)uJ��i3K]VM��$�������8@�r�"0Q�Ed���2x�$�����=�S���������Ť~��	nU�L?r� P����@��6��#'�x�c !K�F-}��-����!k�0̈́+�9�ޝz��7�j�U)�zՆ%N�N����[~��q������u�q
\�G�y��7�o"�w�����,���^�٩D��]9�o��1��1�&��uH��H���xE�V����(��rd�Hxi5���I������Ao�l�z]r��"�O�p�^?������+��z#��Y�|9����{n�·���c�O(C�x!a&�V�+LT�3[�Y�b*̹���w��E��}ȵ|�J���������7V��
 �N�l��sId��5�>��?�X�i������
��o�;����pV�����;�/����\�O������i��܍I����s�/*?��ɡo(��j�Yz|�pi#8�R7+����-y���ퟰ�,Xg6�*�b$m�u?��v�F�r ����y 
�j;���E�n-�iҢ�6-��Tw�t�'ߋ+9SquW�4@>)�C���\�s�@�t��b��ρ����O��X�.6ƁC�e� ��gP/��g����G��x2�3��eU"�{9�����`9j��L+g�1��,�L��B����Lw�^�&|:�;�����b�P1io��
{�4����bk/�BO�. "IH�7�Nd`ɖٙ�2͑�T��u���S�J-Kf�y�*ֱ(PO�Y�Vy��<&��lű���.�j1�9Nr����'��a�Ǟ�Bd�߬�TElЉ��żcʌ�\��`�|�ߖ��#��\���\��BM�6����j��<T�����?���b�D����|$=&6�p�s)5�ǧ�yH����q�!��9,��tB�e	������$����q��KO(��dq1�uz��F��%�}�4߲��� �z��k��`u=��`(�z�\����/?O�#�*�%C:	�(�']ޜO�����Dn�3X �J���5�2��݃�]�$'SXo=��qZ9�O��6��Q#EFv��s���ob�g0{�^�a2�)�HQ���M�,J��S��+�P�!�#\�4ۿW
i��k8��cn����I*�VB^&$�a;���I�1�/m���22b���S�:CoN?:�
>�\pR+l����/���6u7<��Y\1d�X]d�T�ކ:�1ceS�o�������jIZ���X��=�ӯ;�)?a�H�BNsa���H^?�������P��@﷙+x<c{K>
��J�x��#�ױ���+$�
V�q��=%�۷t4�b��؈��@$PI�@��ך�� �� -R.��w���7��}�G�@e���d,��D9�����?��kp��=9C�A����s�s���Z4^�E^�46�s�*���L�L�E}����W�Ғ��{枒6�ȧn�-"��R�Xm|��H�#��X�Ŀd3S̒� ��Ξ���A�fP�d�L	H"��}� +�I�bj����y�|J�R��`q.>&�W^-h-jⱦr��1pM4T�Ro,g�T���=�ʖ��BT���5?!�5g�|zWo���`��a�*�Ǭi<+����89�����l���_e��Y�)�G�f�`��io
@&�����߽���P��3)��ɮ�3X��d�^��r��^��+62y���CEV���#�W�x��&Bؿ���N��Z��,8?���
D�0	�!�����/��8���V����z���q���/q�A�ӊ�'���-��0��HQ%fC�zw�w�YC�������B���R�g��PgX����s�_E��h�k������[�s���Y;�c���uV�Tr>O���G`QoԖF��j�b]SӐ3/�఻y�R����:���0�r	z�l\��~m��<��>:Kv��j+�%v�$k�&�UM�������֑w&�����i���wؒ.�����ty���r$4�G�C���㾓��=��Xl�L�1^�G�wZ"1G =r!����D�eOH�?�K[�$���G4�Ƀ���s;lÂ �oHB��B=��)�>}�cM�Ƞg���ØW���{s�c+�'��Π����zK��	�BO��Cn����`��6�������?��Է��>�Ap�xS�+:ʘ���Ǡ��	�K�����w]�}es���w�z��:��u����7uYz��W}ߒm&���0ռڍW��z�k��������ߕz�d��inܷ�o	��m���#����u}�'��i��O�����L?(�P�a�-�&ς����{�I��?i�|n6ySc\Z�������S�?�s=�J�<Ad�~/��~1�b��~��߷�~���"'1��S7�����rP���
�������j��٬q����\�_�!�vF�S����?N����_d������������ �ت��Σ��O_��oH����KO}��������%m���7�c��v�Z=�٭��<�3�+�2"�<�G�tY�:������`b�u�W_2v���A:>���&'H�����*���у������4��M~�[׍PB��.¿e���E�a8q�*r���HK�g�ݽS�!�M����i:��D�NF��q�u!=�~v��8ۯ�Ʉ��,_M����a�Y��/U�QA	���	t���(���=:��Mf...VVVUU���b��	8���|<^Ohg�>��M�[wm�%�]����O�V(�P\�|��y�iE��Σ)���(�+O2`4��mA��(����]���@����a5Ǚs ��WT�w��I�M��/��׉��$lA��𳎈���o����fH-�:��1K�Nr�~ݼ�ei�A��֯��� / wy�p��ޕ��r�>��9�j����T��g��V�'pz�~AZ�ruu}�����}q�kQI����@Y��jw�K�����*vTf�)
��V_AN��1�O���{�~9�/CX�=ĺ�ws�T�"x�;�/%��)����Ջ���X��7F9�y��GW;�Oא���W����z{�P��?�gDf��o{�P���2�_����T��mo��ǝ�� pf�?�������@NJu�m��.�zZ�Q��_�J���2~Y���ջ�-r:�6��+������-dH] �G��l�;�nm{q��:L Ǣ����ޛ(qcd$�FA�����.U�hޛ'5��,��8�J�3b4�u{�?�M�k�#��~+��Y��3�\G���
2/��T����sqn�O�
G�����9�:Ǩ2˫��zF�>�D��Ռu�������L����՟��{�{���X�|���<u�rz����1Τ~��,����I��,àʓd��9lܓ��=���6�E���<���piϹ{�_b�w���5x=M�Ca>gv��Um
��PM	<�4U��R�Eb���wOi�G��NIh$4���ބ��p����cl-%<�J�§�,�ڸ���hm1 �to��Ɗ�����}�yCl���}>��
;yJ��N�|�7o�X]M2F��6�	;�5�f�q�:\����@^�U9[vQ�.�]o� X3��$0(��/;st�!x�k����TP����Xn^܉��?0�H��u�`J����M�߶giY�*�<�C��qR;d6�w��,���C��y<���\�5ڊt���Q���M���3��ֵ��a�����ߺ�&^^ w#��.��ەۋ���h�F$4�cn�3#0"tâ�ֈ	ʠ���HH#͵�8"L�JtW
`����gg��[��Mă�� �����:���[�D�+�!���`��q���n{.:��EjȮ&3����s+-zFc�<T�^W:���@VMx��F���~���G�k+j8���!"�{az�1�z��<����@6C ���<Z�o
�*���H�yHm��˔=B��vv��=.GM;���c��09��Z�;��%��F_�4��z�����79I��}�tԺeZ�I�uq��I�)z��]�|wV.��ݚ��{���oK������,��.<�U�B^�d/3d�Us��g'ʚ��}�$(��B~O����E�?�9��]��"��0}�i�
\�$ʦ�����n��wd��"n;i�g���9�%ܢ�+�r$��%Էޔ9����؛�z$<y�wT�S� O��`s�"SZH��SE��������yە��f��UL^�Qְ,Z�	�j�Ȋ���j���� /~��/��^6]�?���o஑�>r3�7`6:���<��G��\S����Or�ݱPj�a��Y�,��ƼZ�YW�z��כR��sgt;����z�:$�{u�t]���w� �ʌ�����S|A��kS��Uz�����_�BV?��?VE�B�L�a��u�Lx �Hz�u�w��I.̨�%�A!�����Ե]XNyF����9�배�.`~�"r(:�?Jb��c@�!���#�|�^U�Z8r094��U�>�g�8k^F�m!��>9攟 (���dZj�-^?�%5]+�����O�3@ò����E���so#Q�>n�cܨ7Ҋ-��P�N�TꗰJ��kX��+��ߏ�&W�6?χ�q���ˏ�Lq�Uu��v3�Jkp���hc�P��}V@�JO��_�g�ǳ����.�/������q�?q��&qo�y�q�z�w���>��h�׮�V�+�s����#�&(���5 �T'7Z����6��� q�VU��`��7���,���o�f�̣�b��~���)UY��a��Sٸ��Wr]"-GnUʎŤ����,�c���#�~IZ�����k$��`��0i�9�P@����E;�6��$l�d©f�L��'(�
gjWm��e�ZUz�K���
S�E��rd)��V�j�s�Wg�:��qAJݾ�R���4��4����.#/�\�h��`�_��b���DB���1��b�Y2�zu�WH�5��^��S�N!U�V賩���/YRI;��bU�E%��E�\>���$�����e|6�P�{���d�M'DR-��{R�E�n��4:�a����ʕ���ݭ+�������_i�L�h+l+���@���Z�z�sy���gw��Eܸ�TT��N�ުض]��nh��잃�.����^��.����;�Ua�S�-�s��" *�T��?�?6]V�|]$q]u=�?�V{ʛ���X\QH}�ƙ *���F��ǒy�@y3���v����XƠ�Oщ=ʾ�ǖ��"�#�,6�.;2U{����_ ��C�pKcy��w��Cۺ�)�&#�1�8���ۆ���1��T�w#��~#1��ٓF#��"�X8��vs'�"�;�g��̥γ��J�����' �O����1��_ޫ���HVDV���a��b4����Se�!Ho��Ov����+�t�%0�1��eqQ����M~D���N��"��_�<oa��g
]�Ԃ׮��������y��׻���y���b��$/�R[��h��|(w�$��.�3��䮫��#U�ɑU��D1�i�P,#�؆�S�ݏbAE(�܏�|��t��V<���[��`�(��D��/�D>AeUa��m0�t�����LB��O�X�N� BQ�i�j�3hz�/�޹�{�=�yM��S��:�RQD�&��T��}����cЍ���^��l���-�V���
)F�gϿ�'�����>+fnC���f��,Yk駬�i��FE՛�X����%�c�c���=]�ľ�]
5X9Rv8O�!�������<lfz&)����۠���:���j�9��s���^_���s�?V�W���/��E+)Y��7Fq�k��ʝ�ݴ�Ƈ�Q��?�=Ǭ�n8��9�����/��y�	2(�'��i�\��CZ;r����{{�w��[�RO�Ĭ�>,�&		�z�y�U|��\�����}m% /�'�+Z����|�
��@��I6E���ގ�A���+�z�X����&1_/�@W�g�����U�m<�~�,ɑs������D�2��c�ܙ߈������eߴ��&g'�� J��[��#-p�[8ҿ1K�����B�U�4n����j��^���k���׉�hُ
*/��z�+@M�����V��B�YC����:��`elh��iȵ�X*�٦��n�E<�	?��l�B��@�dtB�h��e��d���o�Q^ڴ�D�)��y,	��iX����7qe��a��S�Oc�
5z,�?lxay�8�w6���2�jX�Ww��^�ގ�&�^� I~�sB]���ٯc~=So]~�:�P�K��}1�:W���l�pd��`=�z�tخ���L�57������ �=�a�ɖs�Q�n~�D�@�����Jo�T�?������Yd�I��R����ɹ���7�4j�j`������£w}T��d�K���w�����vPj��&<1�=^��~ѬO�VPdN�\ڌ��ݱ�]�-��^�q�aN������ƥ�ɜ��#��є#i��??]�}pԽ�D� �#�ٗ�-���.r`�O���39z�͟	-c$�}�|�Q��1&�y�@S�ӕ&!4B��q��d�U�Gβ��n4��td܏�,p�:��ӷa2:�Ļ�c�����(�Jn�w���bI1C��sf��as� ]R�|�.gS�[>��Ȟ�{Д;�I<#��j�W
U(��Q�?[Yp��S�)� �R|�<Ai��{'��s{�+.*�������r����s7?=}T~m�e�w������B�;e����)�l�8XTr2��www=حulז�!'p�E�&�Iu�s_������SAC�&[�C�)�k�ٳN�u]�O��l�'9�Z�󅈯N�%>�+��I:����\-X&wYqգ�}+�ſ5����!c����5607��)�5��-^��6�� �;'g���u)x��v�G�Xr������>'h�l�Cd��X��M��+~u�A�h]�7&�U퓓�����B����1<f��YjOU�%'9�,���(����D\�$x��T6s��Ʌo��e0���y�W�'g� � QA�t�qoV|R�qJ��x!�#2����b��z߳T�໷�[pYø�iba������q_!iL��im˿��E���t�?��s�Lq?����*���|s䶺г��ŷ<BtY�=�Ÿ:l���|�O��;Z�w/1	zN'��{�[F�7���KK+���&/�^�dt���.;�-x�D�xM���M2�o�	�ÊDVTW9V-���&0mx���½
N8�`�:�>&A��,�'Ͳ���o�eHP&4���=v��#���m���I3�"i��L����Ֆ5@��2¬����-�.�3pmm���ICW|4��ݗ�:"�T�J���՗��7�"`��XFb>ia"<N���|; t_``����Y���(í�$cqY�������A�Y+Wa4�m��\/�`
�=�?��1���u���Gp�\k���h�[R�7���I���g��ohu㎳s/�+uծ�)U�v3W�(�JE��趹����Y�*gS�2p���-�4�ĕ����߿{��`��]De	g����0��>*V�X��%>Ϡ�iȀe��m��
� x��6��"tZ�cOO��u����*//�su�$�^��;�뺑��8~Nt��~z�WF�a<�>��տ��妕�AuY��P^��5�TU���q�k��e��/���*N4w��?�����7�t�K��P�U$�H�̴q���8��u�QY����^�޳j��j;���\4D
�G-������T�s����HU�A�! �O��F�A��7wMW�M���~c��vo�޷D����~E65�	֙��q�`b���^ !*=�P�MI� :��iÆh���L�h�		CHtEe�êM����iUU�v�Uw�W�Ď]v���~���9���)�΍���[�R;�K#n����2v��(��_64j�������rzC^fbg.w�!�� �tCiP���ZQY5���)+`N2Iݱ����b̡I1��´�::��k��%�	H�r�4�4=� /ӌ����0���<�m5y��Cj�e�(�x'm�R�̛��^���^�����W��=a�?��~����TP��%���A{�F�'N�D.7�{"բ�������`����@r�~��AVY[�9�U�¦����L�0�	�r�����$��k<��ƽ�݄�u�[���jj��{��%�S�M{��K���.b���(e�m�|�#���?���I#����n`v(��, ���)�����
}��ۙϓMs���jsЃ=R����U�-�f�Z��4W,����m�?�+Z�;�.,|YTS���446�#��ç_19��l'��+i�! �3C���������Y�R/Gj}`�8@\	���a��s.�a��Y�m<���{���T	��{N+�~�5tї(��maG�̭�����2K�fK�}�9����7�V�I�>Ư?t�,؍��"��S�T���B���/�S��8��)r4	�a.ы^Z�O��@�ڞ�#���D�|������(p���6[��ʩ�چ�Yum�5��H���r�*�;�����<Fw�R�����WSWߥ ""z�ݏ8Zfbj��\ �5����8�ҡ���5�6��Nl|�0T���x
@��o��-�an���:2���A{v#���q��ke��8Y"Rx �'xC�6��|��m�#x�kӊ�8�=PAo�����Q>У���o��-����ݪ����o�V�ΜCyth�mmc��E6�p�0�<Д<#IVX�`iY?v&G����z��?�<�@�q�P^��l�c�2�=�cR��>b�z�{������X:�g��iiyz�;L��b+��i��=i����ttd��'�tK
=)U�u��;���d���L���g�{`Y1AA89=���O|���#��M�۔�����1޻�7��y�<n�|����W�S���3��m��l:���f������9�Cm�O��-��������%"���`*���Ҟv&���)#E���kd|�<[({rvFA�["��!�k�\�YSMM�nL��UV�G��徍��Џ͢<��b����(�Cg,)/��M�O�F�,*/qxyyy���JvU�*�A�����q����-+3���D��9 �1y��ruD��p>$�e���VL]`�܏�@,}7��yYY���N��� S�����J����H�O�{�2��}k����Έɞ�C���xvh��}r��q�#F�P�,�/a���r(+{8�{���}�F���6� ��Qb�mKT�Y�K�MMƹ(�|��Ç�����������U�.�����qh�Ye�T��?n�	�9Lf)j&A}�`��|���Z]��q�t\�ωq(B�ƕ!
�����o�����Z��~Y�{�ݹto̟?����l���FN���-҂�g� �1�F]l��<�Mx���|��}c.�[��U�<�	6�;�/�G'=�X>�
�C�ɻ���դ��43N�w����~�Uz��vڂ"�5L���~n����%d���Є�n]�3�=�@{���q�f�[h���4���{��o�vV%�ph�2=����s�5���5����Ф�jkjn�O��<���/`/��/��}/�h�����7K���U��p�q���� 	(cc�޸��in=�ct����$�0�o��	�}dY�wh�<;H���=t�7{?^U��_���Z�CB�x����A�aش�~o��PS�Oym����O31�p�ùbsS(�߭*�z�8��E7xHU�_҈��3�&���s�s������n\g����utx�%�t"�ˎ����Ի����㳟J�����~�����uk�!Ys��/}�k��n	�b�z�Ȼs�Éi��#�2ws��,m���������\��|��`E�©u �����:�UL'�������~q9�B,�Q���X�=U�d�De�D���H聀����ATjRR�>���9����I�7� �Ǎ��_��S�Ygv���������������$|���T��*~ ������gy��H|V&��/]:v��S���m����'&.��[D���������5
9�X�������gk`��6W%�䰝�rqkԷ3a��s=׳��#����␞���!CP�1�k��X�C�O6w4��OhJ�qgg��N��8��`p�^��j&&A��1qE�����j�B3�JT�F�]�=���(��sss}�ɺ��QD����o+�
������dl�x	,����Gd��8E����Y�1��������}p@'���v�0eP�G�`� z�G����+ՠz��'S�<Ғ\9�|'����Of��77��-�mny��	l!� �⾋�ށJf��+� ��F�U���!n���]Dò�}1�2���OSLTŅ��D�!�ɺ��|^j���#��қ�Zذ0t�8�S������fsE���
։ƶtW�zu2��b^Eq�ӧOA�R�C��z�cIL�&�6��h�����Eq����.���H�"///��ʿ�CŖ��?�&��傍v �z`�1υ��$����Ovj*��PW��yW6r�J�}��������z��~�]Z!Coo~H;����������|:�p
���wt�����yȂ���C�:;��䴅oL+�v¿U@!gA! &6quMB%�Q􍫟䍀T���SB�^wS��)9yy(������À�7�\��C��+���&�lo?������e��^��*���(�'����]]�2����9E�(���/6661�#8�Ww���Y��,�X�B���	)��D�O�/5�ʕjc�l||��C����U�I���x�.2�W��1'����-����ǃl��I����N���!�����SW"rX(�3<�S��'�u(�[�&�[�V�.��ڡ�j��v.�v��n�J���e"�PYZ��Л������Ir����4}��{�g����ޙ�=N۶���x�������l�^1�#KK�CBx<o蠁@L)a�\aѹ����H�ٗ�t��aR�b�ݪ_���OO?[�Ä��6�W�ps���\�8X6�"�s���0�tQc�kX�����h��d�GCCcF�>p�}�X��ʖ�_}�j�a;��X���'��Dj�J\�5�O�\v�=�x~�x��Ox²�P�[t����7���|VXv����V#�{<��ދ�����������t���s�N�U�hn0�ڈ��[��6��Mm�5;B�.�s��M��~�����!�q9;�m��������U� ++�I`�����֖!TD�S5d�����&)�%f��+w�6��-~�>���ꩳ������;_v���,<]����h���qNaUko������/S���x}؞�a��oI��u���K�QK���������O'b	E������>�O`���L��}=qssCL
��D�x�1���K�4.�-��#\A�����b�ՓYJ<yuN���n{��W���>��BZ[�
���z}8�i(�z� ���'���ui�oè�["�c|v��x�y�7{�(#�Dx9�3@�����ۂ�<M�G� ��h�N��K�q�6�����aj�y���C��$c<`������Y�>,�b��m�seoE�)�L�jTK!۽��H?bWW�ڼ��`�~�r�����Q��h3'[r���StJ����ǖ;������^?���{dk��wf5��?u**�jU^-6u&B�v2w�e�j�������\Qb��6�%�;ϝ��S0�u���i�F.�k����-.`L��u�X9���I�3�ؙ&��{�@m�bͽ��ڹ�{_k�_G������ڔ��F�M[{o*���EQ� f�ڔ��3fl�Tc�G��w�UEmj�>~9'��|����>�����=7^|��SV�,)���Bc��b{��/�'��Y���qr�h��aų�"
�+��V��=/�7����!���fb
��&����{$7d/N����޾\:�f9�������$�{����C�P�&t:�zw�5%+7��2���q[�U&�(7S)��ط�m�V7��%_��L�>Ѭ�C���@y�Y�"惘�}�׼��?�?��|�V��s�F�E��v���S�g��¾��G�]~V��yђ�]��A)�Y[���q�RY3�gUU�]r���s� �W�t�����_�٠)�,�%0�j�kbg���l*"c�n�|������Ϯ�V0��z4cn8�ǻȅ<wV�~qR�Q����S��+�(Xl��5Nt9��~we7.hp��,�_�4�����X��:w6zk?��`i󌃟?(<&�=��Hw�n�kYZ:��,2�.����|�՞X�¡.��_����ɯ�ݵG�2ʯ�2|�
[\4��Ǹ��t��`9#R	5|�<>A_+eO�ַUB0(iY�^��Ķ�A�s��3�ƌ_�����MQ)���ݹ􌌕�#�j��GVᏧʝ���^�c����v+�3��ٽTn9�=���pW)�>�v�;k�x���ϗ��1���y(�Vh�ZKz��^'��W5�V�Rp��4L�V7�T:�SP��W����~��*�NHwN���F�� R�YFq�G0�Z�]9����Ngr,[�Kߦv��R�0&�I�Ѿ�{�����)��� *�_�)u?�]��I�X��xV�f�s;���wޣ'�X��l��qO�u���B�G��C���G��=:�.�
/�J2��+|,-oɠ�z�����C��������̖߸�عA_.9����8��s�C�7{�U���Wo���� ���A����r
_
�����Kº>	L�P�s�f�0���/'����?�'���m��xR7؆G���4�8�Z~�k����ͩg�꿖0�e�6��2���D/���st�Ҡ��\p�韭q�_K��i!.'׿໨�������]��e���O�j�E��휛("V�{a��� ��H�	<����DC��*�ǜ��4~Ի����T�s�I>�&�yf����C	\���!�x^@�wNdCR�%D�����kO,k߮�R��Џ��.ܹZ�Cb`�.��~�{�6�����L�"��_��Mm�J<h���B{V㔳N�gl�WæC�j]�f�j�b##��j�����v��a�@�8�*��\O~^���Kk.7��T0h��f��T��p�b�I�x��1��?�_=2i�!I�&a��D�Yd��#^���Om~�"����Vt�B v+���[d�b僙��h�$ 5��-n��[Ӂ��7�wH�}3;��???�4?R��R6/@Y�!�{��1���ȼ΍e������K������Ԗέ-Gl��o��/뻹�H��۸x�'[5�)L�,�|/ڒ=�
<*/�\
�C��'^MV)��ğ@��]u�|��_��W�0���f�u�E��&��f�-�R�p�V!���N��=�L��i�s�՚ue�~�m�2��d�����~Y�/���SW�K��|�i��]m�E�KΪ�[��8?R��"gS̹������&r�]dd}o�q�I�2�� ���,�K�-1�'~��/V��<�6;�ϵn� ����6C}����l7�<�e�J��Z�$�9P}�;�"*�싍�U87���?�+�MϜ.��vs��z�;���Ɓ�\�-�O��tafY��);
J	z�{)�QC���1�(jF1�>�G�k��N.�b&���y�0勨9��Z�Yja�t-T ޣ���y#�5��2���3�}@B A�+�����M4��6�MCHŔ��AA+�B4[8}�@☴�4�Ρ�Ck-����t6���[
#�;�'qi�=h��b>�I�γwJ�*%�xpo�u���Y;=�k^��K3v�t
�O`��"B8(L�-~�@s������m`�7/�a�f�):�ࣲ֞M����ͽ�B�T�a.�/�@�����,n�@�q�*t�33Uz�
��朕rZ���ٷX,ȥ���&{U�6��G�i�q��X@_���\>9$��?��ťxB���a��{7Y��X�Bww����F�/Ό%l��e���U�|wv�:�!!���dX���M��]��l��~]
�:����NuN�gX���I�_���hS��0�"&|#�T�Oּ�����P۲|�t]_*\��wZo���XOU�<G/��U.m��� X�<%&%e?�e��T?O������j�-5��Ǐ��X{ ������ֿY)�#����{���. �>o��A핗ޅ�t�3[*[��U�\~�8�RtT@㠠̾�>�n���>��$۴'[s��������#�o@FJ�EA>���ڥ/B����D�D<V#�.J�e<�c�;�'��J��U�OC#��L.�����bU��яE�Y0�Ա���<t������Q�ȱB&���z��(pK�Qrr/YR���%O���M�7�9��_/9i�:u�Cs�r��Fts�&���t{�Cd@E2

��wS5���� ��!�V��U22�%�|¬����쀴!��:�ک������'�v�6V�ib�?6m���u��S�2�Iw��bG��%j�prW��"푠ZA��n�na����ls��*�鞑Q��o�[h�g��������[�p��zSޱ'rI���ƿ��%g�vօ�����leg�?�V�F�*�sS�Zn%o��2���P���.و:Xƹ�~��n�ݿ�H���Iβ"�sA��<�}oU�����o-�6�k�E
�7���q�u?^��w{��m=j�15���5M!cT��	l�n��G������)�N��Ǩ��٣�.&�߶��\>)<�?5��Kb���͹*g��Bq��ɬ�N�_��Z�W��ZX�\s�j�-=J�(��&{b�pr_aa��K��h��x� ��H��du�ݦ��Ĩ_�؆�>�>x����|�D�R�'Q�@�0D^R�P��� �\�ؽmC�Z����`�˯%�\���Z����>��&11�������x��8uNɎQ� ��ɨD"�zA�C&'<^����4�eO�|o�D�Vɑd����~����8=�tw����:1cB��yu�:4�g5�$�l�J�m�qM|"��j�K�iN��b<�
ٝz!۔8����*�L�3�򿑸�M�a���\_���Ѿhq9nx
2'&S�7&AIj���o9L����7N�~pt�<w�8����S��&~�~�!�	3x�YF債���=U�HM&Y���SL�H�_-�'j�ܻ�o���y3NT�J-l��2�$}����^7b����� ��ͤIA���չ*k�2u��n9��O�������v^r~��_<��CQK���o�{�Y3x�e,�ϝ���Mc���9� 7�YN���E�T�ozBKN�<�E�n�h�i*����3��:8>l�w���O_�Nw�dbGwXW\V�ꔡ_��|:��'5��u��g�k�)�݅L��=�=��G$�I��~�ы� Y;;����u[�rБ�1¢�mă��Omw+�����Ek����s�U'�,.����3f�{�a�ta�uxA��(�t�0'���	�a�cI&M~K��>�'3諫t���j��fi;���	{p#�֪[�oqf`��(I��<�ϥ�;/5��֒�LE�oe������l���D�	bj�p=�=6���7ޣK����΂���544�r���U'`�����7x��y!��ɫ�E�
�c&��l�/��Y��.��Cb� B#��ZJ6܊��m�,(�˕4b�����9Pǔ����E�6r�#�z�V)q|ɇ9�P��FR/�6I��k�XdV��Ve�Ly��ߖ�kp?��1,᭨'%�%{��e,]�$�vm���r�x������iw�ʖ�8cW�W/O����v>q;�;�$�n�F��P<١�&M������?o���k�{
���>�M�% 3 C���Aoݏ砶��#����N���6��Scfk�/�	sLi�f�>J��-J}ޤ�9Y�gCf�7�;���$��\w�*n�t̵opej�Fv����5���\ﺋ����L���-b���N��(ڄ���g.bXoU�����p̺�IX���j�u�k5��p�������W�s��;ƫzb���D��┖	���6#��͡(	3	�Rҟ�,z�'��W.$�[%J�����>��I@-�J�z���������&�|� $<3�t�e�!yέv�~����q'ɛ%��л������ـB�F�¡�f����x��gZ��lm.�c�iҴc�W�צ�
�UY�u�3}e�v�����y����+ƍo�d��嶨TY�-�)+`I��f�r�M"�M�	�j�9��x��J)s�ˎ����yhmy�A��F�z��}�����F�s�S���b&�2�ۣ�Ķ���6�C��z�GS��0��c��������H�ȳoGe�r�Zb$��.��o�~$/?�p�?��_SY)*�}	W*�1��"r}�#����"�������^O�Z�F �c�hƬ7,g�;�뷚OR�]�zp����W��]o�����΂9���~�X�'�����ۥ{HϨ��Y��+NNN�(�B�B��]<���`,#�!h��Ae+R]����`%�1^��GC�d�ippp�^��_M��i_��^4ZqC8��0�q`�����*q��,!.(� �0��m���TE�O�Cz�tBfb�������\Qa��y$aE���5�MLu��?k^��x����d��6%�r;+װpз��ak���Bg�݇�O�n�r��`ҿz���ެݫ�(�"��Sݜ�>���W�Sϙ�2 ���=yv���0Q��k�zgɹ�!�r���6�Nذl�� �r��B)fn��`P^�F?��|H�+�nէ���1d��1&��S��ē�{c��'��b�ܾ/J�L�]���.��Xצ��s	%
�VA�����^��SvE1����L�UW��-̏�G�^}<�o�#�9��\bY6?^O~�*Yp;���$�5�:�7��6y�[�9^��u�q��G|YR0uh����g�]K��(�뉯π����ߵ� )���V�>k�:�W}k�W� E�HZ��ݣ�ލ�-W�xaR���}�;>�[�[�U+|��8u��a���$�o�:�����DJi�:�e��v�L�/��'�*���qn�K���O�b�4��*>�հ�''���IBH�u<�Ue���A�T��7�X�2Kc�sJL�,�ѻ���Y��Y��e"����YR���:B,�].�*�p��n�лي��Lo����ɫ�6�W�Z���N�̲��#E���%莯����l��A�A�nM����v��(FLr�N�d�}�67��@'�����K���ʂ���۠E�E~�]y"2�"1���ms{>G>��zQ<<c��bv�\���c�?3��-��n��UGKm�lן-ݛ�[/[Wk��cn��>-�Hᑱ1q�X}��aM��UUM��M�DnpZv6�T��A$�Fv��r�͵ ��y1]5��[�W�!�����Ӟ���*)a��~�<�t�͈�c]w\�XX#�Q����ԉ�"�+r0rV�E�~=>E6��>.)v=�b��]��III�&˱Є͸H�����K2��8�>�͇�<����rb�I@��P���o��\U�6ט.k��ֈ�����w��smnGJ܋���KwO�ȟI��ڜ��nƁa�zSW�\K<�����9��O�y]𛂶 �-�Smd7��/ݵT�:5��D�~�����K8��A,�b��VhK��Y��LW�i����e�y�W�F�������<�I/���/r���������9b�]|퐪-��0V~��j7��1=� ..�b<r�8�$G4j�={m��Tn��1ɰ���x�3�5Ԉ�핛��Q�H�n�W̲�~�W[��1&��"�#�I�9�1P�:do޵V�KW|Ǆ$�=�<;*!����ՙl�<�P$��*YE��� ��U
*�hBI�U$V�E��c�]�Ns�R����<�Q;e�`������#�}z��9���.����~1���'��  �9_�|s#���v^G��h;�r��l1��䑗&7�z$ ��;�Ȳ����������{t��b��E��ډ�����#�-w�W�fo~؊�51��t�Kj릧T�WT�rU9��Q��*��R��=��4�����q���.����hK����:~��6��M��11*O^8Ì;"�\2���w~03)v������Y�#2VV}�WZ�w��C(O0L�t*"�d�4S���6��48�I�Uqc��2T7RGs���W��;z{K�^����mF�	��P�Q��r�q�Et<�.��p	}��Nl<:be���E<��߭��i��ScXm��xğ<����������B3�*׭b�c���#;Gµ����ZP}���b�	�|�,yi�P���Oa��Pc�������������@�+���Y�^��{��W/S{��PK   ���W��W��: �: /   images/5eb2d398-7f6d-40aa-a255-437b4468b1bb.png 8@ǿ�PNG

   IHDR   �   �   Z�Pe   sRGB ���   gAMA  ���a   	pHYs  �  ��o�d  ��IDATx^��w���YЋ~Gyۯζ��%;�Nod����bC="�
rE�1(�EG�"
� � �QD	��fHH٩;�.��Y�-��?�;�^{��x����Xs���-�<�3�>D�1��"@�Do�Rq���<�ȣ�v�=�������J!o����摋�����+�B�^���s��	�M�~�#��� Ā�!�KcD�g1���"BD"�d��9{���z��D "BH@�|���SC@J��:~���~��-w�{?�w�'�#�Ǉ���'������wr�w��_�u(�y�cC?��ol���I����P,f���S������O�{���*ϖ��YLHJ����?�s��_�ϼ�������{@ ��^��������]@�}�~��S�=!zBG�����{����?���u��)|!�WJ����(8s�m�`��m;B�x���=�u�	��|���_���>�j�z
���d����Tp���ϵ_�ޥ_�`��6~�c����p��%Ξ=��Z�~����!^���2��n��������B�O~�ӏ��.�<o����z��˿�j��H��O������{���iۺ��}/��|죟�m:���gx況����3;v���u-��H�!�;蓟�l�F?G��r;ƴ���п�����؞���gjO7~�Y���I����S���|>M��eJk-:����Ci������@Bț���"d�ͅ$�r�,GJ�b��n���>|ύ���|jb>��k[~�o�m����?x��� �<�B<�z��4��ii���/�$O�v��i�|�v�X����8��C��1�}����>O7���1��/��B��:?��o~�ux�8�@���q<�����8�
n���_� B� Zk
�)�k�X��7�~�;<��8���<�q�������
�IΤk;vvw��m�ق��	����B��Kk%�Z��`���s�-_B�G���q��U����e�x<@g�% 
��/���?>/������w��FL��h-D���qqI>����8�.d��^��DV���r���ȟ<�eI��C8c)�)����oģx�Nӎ�w�Y��w��`�s�����u�g}�������nD�3k[�<C
��ӿ��S��>+tm���.Jh��H:����^�9|r��
n��՞n����y�����BH�#�`��d]�X�q��'�6�g�M@ #h����Z��Ez�M��&����p��:��cڮùd0�1���9x2R?3$~�n:��*%�d�wc��=5<�O�nx�s��rI�2�^=�>KO���{�3��4e�Q��u�Y���X���>�d�|��=�|����&Λ���>�B�C�e�͘��b�)g�1\G��DBg�G��"�QB=k�xZ�D��VU��]gq.�!�<O���	��.:+0�����L3vs������Zvvv��C)u�S�3�σ�=	f3ں�i;����؏V�(ʦ���ߛ�|7_�jO7_ws{q�L�7S����ԉ��}�$D�p��c\<����]�"��y��|��5p�$�a�}�24*fd�&��NI�:�͟�]���'��<Zk���m��� �-�Ck��5I��!��̛ۍp}qS�h�("U^%�@��
R�n~�S�'�7@"!x���\:w�a�F������gȾ�F�us;[��ݝ]�u�Ε��bB�D��(� ;�S���<ӵO7�{s{q���	�ャi�5�~aC�y��A��C]���aC�H!PJ���9�R�� �f1��"D�։@�
gl��'��̓��y��Bb��)�(�
�Z�HD�~ȟ7��b�*"MӠ��XC��d�B��7�'�Y��3�f�c�`� k-��B/���y ����c����>�8/�����Y�H%���`�w�zNC��	>��
7�2ƈT
%]�]'~,������:�=?x|�(�ɳ�"�L���X����Zȧ��=����Jb�x�6����s>�0'�b��C��s���������iWRF�q�|<��)���f�}q�~�8��;O���Ei�xo���ތx���hb�I���c$��ݽ�|�e$O�Bo�k6����"�Q��?w���GJE�)Z�Ҷ-��^Я@�x�Ȳ�7��<�7�}�ןb�8��ʜ��8�������-2������J)t�$���s?"�]�@R
���="&BR"�z�do�'���T2Yc麖��Y��Ig�w�g���{�뮃H�y��)%��u��6W��b�B�֨��q7��v�dYƠ��3�Z={*�} �ȍ�FxJ��������<1&��u�󆨋g�_-�R��D��@DI����O �|��Z�"c�8@��X� CH�����Y�ߍc:��{�hU=��ӽ�s�+�>�(��)u���{{����;�Tky뭷p��-�E�ֺ�y7<���7��7���&Λz�?��1��s��a�U��S��!�2荟ǧ	��}��)TPHA�+�Xӥ��h0��|����	�c�3��Q0F���Z��δ��K��<�wq�#z �r��yL�?�	/�})�5�4"�Y�R��������8k�x�h�_wu�[��Oxc"�C�ؓ�(]�8�	)�Z�X�PJRUD|�x�A�������w�؇���k�����g{��/�k�{B�I$,��<ט^|c�)�)Ɣq����H���Xc�ɋ�ݽ]��L>��C�E
	Q�u�988x��{~&�q�0ס_3)����똾{:���O~�!�H��`ȴ����D���s�'!�6�p�b>'Skkk�g�&��n�����4�:\��S��p�x�v�4�����-���B��$ךh�9�u)#F	�ֽA����C7#�S�+�A�)@
I�e�t<&�֚K/����􄧄���q=�M��F�>�������AJ���tp�J���!�{n�?}?%ܸ~1F��;K5���ޏ�	���<�l�f�y:b�������5�}P 7��譶�����'N����KbH��"(I�3����ۡi��>��D1��Y�c�e�\"��C���07 ݳ~G)�7�V�
�s�OVo�OU{j�y�|������y�Z�t���=�8�?�YGU�L�S��I�����W��\��It�S�A�ڦ��C�ϖ8I�J��1b��}�St���b0���K۶�p�޸���#D/:w�loӵ"�d2����i<=Ę�O7F$=��wR&K�����ѥ�����Ͻ�HV����-�@�5� ���wq������w��;��Z�钏����}��;�=` G ���Zb������
@�4y���@�F<w��_n�j;�,$B�o!�tap2�	�R���,J��8<Q9��Q.Y$�� �~ Bh�X,��$Dׇ|y��lh��;�����41�dŐi9��Q>��O��*�H��'"�o����R#�	A!���`���q�����7�� ��@K�p<� �"�� l�/�k�݌��:���(#����Ղx��C?т7D���ۏ?�p���bGS��c���Ap�8|�i}�ot=�Їv"���>��-��y�cd`�\�%�� ����x�Hk��&Bx�o��O�ӣ\x\�z<=D�'���z}L��F=���tH	�HTҺ:���u�s
@"�}D'H$2J�1��� !QA�}K���R�%�&I"���ƞ�FS�"d ʐB�dLT%���+t��Q1�rBӐ�4h#Jh$��5B
��U�Io<WK{LO��
!r�P)Ah2U����GDϖ��<����0߻��M[�gi��E����Ϩ)���H�(�b�Te�`0DKE�4�|�i�p�D�����D���$�{��:���'���������4D�A$WQ�}��]_#A@���A��i4���u���f�l� #Q�Ħ��t�~9�HB�H���
!�ei��hY��BL�}�R��^H�)�($2�~qt���z�	B�Їw\gLJ��/��ˈ�O�'��H}�2}2
TD!�R����h �Q<J��1CƢǗ4������wD�7��b�tx��=bzE�'"�����I���ճ�D,�D�8�	7�	�*���)p���u��v���\�!ڈp92�J�'81��g��xX�K>�{;�#�J�d�d+?B4�m	�W=w�~][���Bp��,QG$�`b��8��xO���-����5-�x6F��`J��G"��<�
%:��.a��:|Q�xAw�7)I�r2U�� ����D��<��%�o�_dBp'����x|�$1��bA0�51ZD.��"!E-���T"��+�d�'�#�i� ����Le�b:�5��D�T�'����*=�zK�?d� !�#/=���oVD"G���KGNB�i|����G�߫%H�1I���&��<���v^
�H8�?�:cQ�h2��\ ��� �"Oy���v�B�~!�D2(�ӏ7�Q^#����
��d`�D zZ�ܗ��FZV�ø�ϲ�%>jD,p�@�k$��CI���z��O�zZB@�2�S�i�;���&D�(Y�:�d�N3oY�/ɫ1Nl��+�N�m5�j� GD��"Pj�2+��tƱ��Ǫn)�6փ�`�ʐ:�h���9arL�O�훓Oq�?������Vd��6C���N�lOᒐt�^%�}��Ĕ� +"Ax��,]G'�H�)"=Y��q��)&$���t���1�$���Z��β�?c�;�DGcVx���q0����	簥ϒ
�H�:"��+��<�$/�1RbX�H׳�h48�`�0��)�B���P�!B�*�Du�ջ@��_ 24��"�M�$(d �}�}��"��D�a�@���(��)������F)#J��&"^���X5�[ҭ�E�¬о�}��5ĆI�d�Q*�� � *8�D@K����P#c�,5��f.=�v�w3r�A���2K��-B�,�?�G�^�B�$��NrfrN�`�6x�w���Ȋ����p �!dV���*���:��=�GtdёE���[*g�Hijr�����P�R������5�h\$i�$l��%�����s���;2�P�m,��za
�
�
�A����'��BG���bdH8,�����;��m�'}�¼�܅d[1�c�~�Zu�)M��`�-2$�A����Q�F��S�ZthоN8:��Dvd�B�6M�!�^#ڈ�@[��e�k�M�j�#7��
�N"�l��B4�=��Dl�u}�����N�]1s�m�N��{�;t���X�8k:��C�D�2���q1�j�'�^�$��b|�+�������z!¥+��O�$��H>Z�/��?������+R� �*a�Ƶ�&�� 7A4��xt���{=4���;?�/��ފJ�׾�����C�։m�k��v��~뭼��/e���P�z�)�I?I����>��q��E~�������Q^���x���#���5>���3���dckd����I��z�*}��`A! �i�| ���X-V��?�s��r�H^���c_��R7�qu��[�H��b��C&q8�=��Ğ���H�������[�� ��q���[��;�:��["o��Ý3x�z��AGC���R+���Pu�����.^����_�ʅ+L�ȷ=�J�w�1r9zth���_���
J?C쳘�m%DH�\���!Ð���'H	��>�kQ�~s�	?}Jb�"CDEV�t���!=�~�J!2�`�F1e����� ��J"�w�I�v���.��}+�-���Pe�"*:(Ek:|��� �-�ud!����8�h� �Sj��Q#=R�@�"n�i�UJ�K��t�զ�[�Z~��9�r�`��޶ɗ=�6�L2V�!`����=̷�2��R`��Y7��� :/�V�Hc!�����5>]e�<��+OLȜ�yG9"������(oAz��cyƝ��"j���+L�@�d��.	I!�)�6���9ǩ�e}� /}�^������I��#�;W�7����E�z�Ɵ��\:����2�����&6@N�G,� ���.9�E>83�n�ۖ/;6�EC��|�K���7~�M|���Os�C�a���L�c$�@a�Y��<���I�,�mI�ů�W?��:�bz��^�p߉M^��������W��`��9�[~�O��@ft1w�P6 �� 8G���\�/�����]�?|��\����c�n�Ɖؠ�WYW��9������eD�@�)bO��(4!t���P�T��aA�:�ՅZ����t֒����t*Y%u+A�<��v��tX��S���-����(�YV�y�w��@�~�m��/Qo����F� �X��=�7�k��d�cc�E�7㫏�����6vϱ�s���%��`r�����?��|N~�4�Kg�}��/q��9N^=��+�o?�x�1���Rn�c8�J����EƳKT���]a�<�xq���2��9���{W`�*K����c���n?gs���O��4��8�K1��(Ev���G����[��ｙ�ΜQ��`o������0Y,����~Þ��n� �_:E�-i���Y��]�1���L�����D]��w��^�j���?�N��`�
�C�J㨬@��+��T[rvt;�V�[��w�I��#��8�L�"n3Q��hq�x�Q����f��1�`\KF�a$#���/�bI�CͰ�cU�84�LY�hn��Ӱ��c�U_�[���������کG����]i�()�����\�#����UG��#W���IZN��.8V�[['>���W})۫]�{� 6oGV�����JiJ�P.��&S��{��`�����2>�
>yz[W�]m�
r�:˴�jE&%�R�,PhI�Zdh��d��
-Z�hQ�eY>Dg#*5��9J� �@7�*B���1�݆2����}1������x�KGnAl�9uV3Ѡ-����Vt�)TA3b> ����B��n�+1��v��p�]�i�F�ǖ�(._��ڠ�-��)�,��[^cOd�n���	>�u7N9=���d��b�~��%�%��32y�*�c(�`X� 4�����PGѭ(�����22�3ʖ
��ӋK�-z��dg������jH'a���Պ��2�tKD�u��E��x���hu@��e���K�_��%���]@5`W�Ҕ�3��?�z3c]E8��Wg/�Q ��k�=�
�X����*Y�m�1��ӎd�]w�1�-�`��#_ �AG�Z�n�kvp�+h;G����.�0��9�b��\H.6%��\�vi%�-e��v0�f�ʯ��%E7G����]���]D�Op�s�hv�f���I�i�t�tW�����Z�n�$��`���r��g��� ���>�@����4��̣h���W��)����j�Y$2'���}�s|��k������3�	��]"tW	~�n���Bh/�˰<�e��"���YH�=0�4��O�c|l�E�������~�;���p�w�-n����_�a���p���I���|��x8L��PwЮ�9 ��6��ɀ'�ZR1Y*%����	�5`f���ػ��=�.�ry�a��kG�!��˹���2/�޿�+����G��g�:����7����\^����*�4͂f�t�5�.b�˸f��o�fq���η�����_$�Β�E�96*�B2��
I[�L�9��f4Q��0f���-/b�m��7sb��[^�73���j�C�g�a�����[�Q��ְ�3#Z�]�5"V�0��!t4�p�5l�G����%�?O�h�c��񈝶�%j4���"�d�W0��Ѿ�%��h�{�.~��贤*2���\�k�Ѷ��⊸��;��b�4��<"8�.�)�J�1V:�_
r�ɋ���g�(��wq�}hHۂ��̒�^��5�̠�	�2�7t���6F�A!]�m:Кa��"h�Π���+�|�%�`�L;�{KG�.���K^a��Y�v�	3��C0DS�L�l �!��6��t��`�0Ɇ�^�n;L��s�t���c��c󋜻����^���������W����w=��-w3?�Vǟ���Ws��������/�}N��������K��ۧ�p�Iy�}t�� �Fy�@�#\�:.�ϱV�v`���'9"��{��y���1��+?B�����]_��֗�|�k1_��|�_b�;�����y��� �5_õ��Z-Lf08z�lr4�hǢ��EQ*����dg�i�X-��+�Fk�ʌ6t\�K�J�_���v���-�	�s��_�=XB�8`�-B@u��%�옴��X��{��8`�c������>�44�£;�3��%�k�,��CU�e�@���u�tH�B�q�+6*�
� Mۢ���֡�fw�*��.BGt!i�u-��]�5�b	�V� 6lFO�:�?�v3Vj�=b0�< ��LB]ϐ�Ѷ5��pV�Gϗ�y3G��V�`u���udB1Z��44��]G�5��bێ��L���e�L�/S��B�!u���]���j�$*L��Y�:Xu�td�1X%C��@��yR�X�<��b��c�s����&٥���������/gw��vc�	A��$��<(|�S已�������������x̴�V��p�k�~��,�B�p��OEu�(�
��ˌ���'�� ���^������l~�?�����-�t�F��q��{ɂzy@���u�|w��˭�'X���t�:�._�ۃzwA�(f�vԳ�n!(��j�$�@w�=m�p�%�4^c�^�#�Pxd��)�
؋�E$jX��P��-ȹ�FQ�S�0�E��G;w��#�D�;�s��"J��)��,!���dm.� V��Nqi0�dS������!�c�!�[_`�A�3��f@YA4����D8�O�py��ג�0R-s�<.�M��?ʑɐG�]=F4�Vk��c���/��
eA,t�A�H���9�=Vֳ�l��5�%���P[���JX>����Yߵ�^�fmc��s��[\Et�m�hW
j����lI0��J�� �U�r���G�\eA�.	D��B��u��Z�pF&�r}�����
b'�&?<@h@/F�f5�	E����Ky���'����hu/��C$c`�[���8��3��;ͤr�$�f�z���y����8w�����s�;
+�^��9��q��� *z9BE\A������n���?����
!�T!2��Q���Co������y/��P��}��3:Ax�q����d/52�ه� ����c�� � ���-��8���Za�$����Y�2��Ҷ��ej56_$n(;pv�8fցl�:�=�Y�+��b�m��;�>��
��0�9�������<��%�WtM��9d��C�!�1��K�B�lI7_��[�0�l��oց�P[h��!�5��;���dڦ��֒-�p���ł�C��)�G2��_r����"!H��,�'&���.�B�/x�^bc�g�,��(�s$�\��I���Q�f�[[-�� k#X��P�%�j��Kߢ��p��$�WBa�g�0�W��!�	E�r�M!���Q����4]��ץ����8� ��� MrA�]����W�����g���_�*J�(2�&�g��7��Ͻ��������-����-���z~�_~/����`u�C�-Yhh]d;z����x�_�������&[���.E��;'�"@ z���ܖT�8{�f��]߇�گ��a��1i�y�O�m~�o���������ߟ��ٟ�}������-����b�\pl4&��&cx��q�_�싿�Z$7�]�(��Ddq����C�B=Vm�~�&}��!k �tT�X|�2��h"8��$���8A��"�;�$�x���7���	����(�YE�2�)�Fuf��].>�xe�2�wd%:�4}a!8��I��R!�%$!ˡs����TV���� O-?��FJ���Z�%qe�Z�[Ȼ�n,�ט��o�;Y�$빠�"��ِ�]��%��A*BH��Bb0����m'�>�'[G
�߻������f3H�����qY+���rb(1
Ԫ�.����}`%�k<'I����e�bBW��/�e�j��o-y��Tr�z��M^AbćIKJ)��R蠈Hy�fOA��%8�mz��?�7)��i� �U���}���_�Λ��ՙ7sϋ^Η���_�����_�eԟ�9����͟�>z�/��JedbE����=�.��� �\tw1�v{�o�ϓX����G(��\mٗG���?L�/&VcN���>��������o��<���#�^��7||�/��?�=���(5��O<��w�
G��h��Z1�>�26��`�0�a�C�w@3[�ɴ������y�7��i��kAВ�u�=Y�[�`68�����Bz�!"M�Y�|ˎ�K�~���rq���{���E|P�C��Tݡ�*���*f��rw�uh]�[��AQ ˎ�Y���,�p�#�7��@��9F����D�V@+!�&"΂�!I^�X�DC��(���� i<�%�g"��2�0�eJ����#(I���G��$Y1LA�}0�iSdS�cDH��tM��""ŗH�"^�L��]�ۼ�6�����x�:�l�{�N�'�-a`-@� ������;��������[���^-p�@yO�4Jx�fI��"�Js#�L�2�R"z�C*�i�?�L��"�Е��f�/y �5�}=��9�h���o}����/�v�������ۇx���'����۾�{x�_�����e�y�>�O��ϼ�W	*cT(�L��5F�g9��.'��dk��K*�>6�D��[�,	Ns�;`�䮯�6|y�2*ʃS��G���J�t^��y��������Op�}���o�E_�M|�w���~�w����{~�[���cz�������5�eQ��Z:�\)�=��CƤw���,��|&�|������m�屓�s���٭�p7@�H�fi3�3xl��7}�(��7�q����H~o�s�(7�0��mh�H�PD�ΥpGU�2����,*��o���X6"�p��
�t���g:Bעoj�fI�,U��)�K�0� u�հ�i�_�dH�W��$�Z� M,�^PX����8�㙢��bT�����.���L�� �dBڍ��6�t&����Ev�79{ �����>�i~�������\.�2�IU�3�I�r.}	gn���y����@�Ż�pi?����@U��=��O�r�
�]��> |��ցm|b�-8q6 -�]�K{������q�B�:�/������G~�����W%��\�O���zz��/�z���_�%����W8��?��@A�!�p��^��Xi2�	��,���I�r8��B�p��<�^�EA�`4����-���ϗ����5����PB^@.��ʊ�r⋿�?�]�O�*�oJ"W��i��b��5��g�t��d� e>�,W�I�:ȞsG��=�b%r>�=����2��:g��d~�� �	d�`B#
.K�X��o��2��3a�rz�8=��C���`]��5�����'Ĉ�
Z���+�U�2�h��̸�J�-$�2�1R \ ���,���#+�ת���Nҙ�:&�p'�簊03+���4\�pJ��;���`�:/6RYM�'$!,�s�W3��
z�B�2�8)}��axr���!!{�H�.BA5ޤc�Z;��ф�:�G���Ę����Ę����5v��|��7��ߜ���>t��.=�������n�z��;��0(
|�T���҉��!��p�V��^p�� m�\2�=��?�:B�@�����w��
^��o!��Q�Q!EApB��B��[yɷ�E��~����w�<��N�\�5�y�_d� )�	�ύ;�<L�~DgQd�-�{����]��P��ӟa�Ϳ��+rϷ�(k_��,�R.�2D���t�B�[��ʯ�:N�fw���Nމ��4��1ã��B%4]c�!�F�G̔���3�4��|��`�+�.��5cxGhy(�\�PXz�������C+����YL��*ֈ�B��:�W}����!�Ze�,c��q=?O��Y�e�C�����P4���p:������R;W��'�O=�AgاdQn��>���vFw���}7a���n�z�s��c�z.���?x!���N_���\8�<N��SG�ˣ�)�+�] 8�ReǪ^ �����iPd�v�L2�yh=4m�=Rq2�N��$�K���HhWe^@��L7�SU|ZO8�r\6�[(=�;�WL�4��A/���<J�;z=]�Eŉ:C8K��1�����"�PdD.p6�wK!�t�2HJ8A���m�o,*�L�����R,d��O|����5/���à�Ӈ�x�qV��z���6Z�&���8w�����7�-�b@Q�^�_����i:���a�R��[D:�%�~����{��܌av��}���r����9_�gh���Y��	
bTh�Γ9������'�̙��I�)��w?��u�1�zI1��nV�.��&�ɺ>�LKŚ((�t噘��((Ąu�Α;�9WgW�VD��-��))��+ȃg�c&���%��@vCD�Y��B�C�ɈS��riw�
L�����L��B*�KHC$X�H̋g�K���yק���{��W�up��M��-k��-����͗�����㫎_�׎�[Gy��o:r?�u;?�~��Y?�On��W�[�/��Vu'�Vl�NYp�������X�����ԋ��)�$+'�.���R����>'��z����RAq�v3Fa�(:��%�vA�$1bh�>��Mk�]�����2�����4�3L��;5D�RtΣ2Ͳ�FQ�Rگ���\�@��AdV���f+�G�)���FJDr�m��%X%�ö{\�������AT��E�m���mk�Y!]��5:�)����l~ӏR�W�Br�&�罜�Ŝv�I�Oq��zM?�n�U���w�p�h��[^��4��m|��E�אޒǚ�� }��")�A�W��A��;G����V5s
��aqhq��J�v!��6"�}o���.H���BR�.���6��M�B�O��D56�<�\�R%Ad,��"�IAn�.�~�T%e�����.@P���B��Tc(�$�8k�1`�^$W)���T�.X>��w!P�@�3LU�0�=c�����{���V����±Bs�Jõ0d�7ّk\ۂO�r.�{aĥe�c^��8�섊>/ЅNVY-qQ�,�K�Fc�Հ���}^7Na\�YJ/u��L� �(2к�t�T�)�t����X�'�\(��0����aO���N��V��z̰Xc�@:��0��jX"
M�Ȋ
�g8!�$�F�$�V��b+�uˇT�A����0�I@S��j�������탫l>�.�����t1�F���ǎ.LPؠ�!��.9�����˸��Q�E�u����2_��K!����DI�h".�Ѣ��[r���/��<)�ΐE�Q x�.��Q�Jŵ�HӰ�����|����W�*���K�~Gʊ�
�&��kۋ�J��)���!W�8�,QBw���L�=e��;ρȩ�5t̓R��XVx�U:�G�"�Q�)�B�Y� �J�@��9��|�x���r�G�>A�
���DNAE1���cUI=S*�r�r2Fɂ�2<r�[��<�nG��k�b�A��0#�[��� �����\g8o�J�dA',�Vd�yCpIO�5DrD���S�.�1b]�1`]�D0��uq$Ȅ�FXDV��T���"��Nh�H~�:�TI��T�m��5Eעm�)��	��4��" �48��9z�;4^��ZC�}����'U�.`0cWIR 'w�V�:cw6#?v4�cz�B�H�F"`�I�n�8.@�A0>z?}�֡t��g�!ӣ'�T�>ѤP���{��6��O1ƢU�Մv�Y� ?�b��%>Ę����kp�W\M���]��e�[��(Qk�[��+�cX�V��EBp��#$hK�\�x0�����kR2�%s�1��j����qŞ(�3VB��%r�^��rv�Mَc��&W��9+V���"+VX?#k.2�*��8�ұ}�}LV`Qd)w�y2�L��`����#��Zi\�5��F=�n���X7��F�rDy�ɖ��a��t`�-^�(Q���n�K�P+�z�x���&Pـ�`� ��8?E���	l���DJM*�"4Z���(��E	E1DfI�Q}v�y_�DbbF''�b�U��*�0�6�b�*b(����hk��)W�Ɇ�>(�]��J��d�?"���q�R�cz����$Q<��&���tĬ/4�S�%ES�#Ʌ�^��P/�$�n��J�jVPڈv��Gr�D�9�7t�b�C����ɻl$��9P�G�Z%����#�=���ɟNﲒɼ$m���.��E�|��9J��)�c����%�%�w	YH������A��4%3��D���?��B�M����r��$N�-&�T��`(h���Е��jF֔1�vJ�� �%7��1��:m��I�0�p�r�Hŧ768s�+�x�UlK�{����2�-'�d� �0�'h?dUj��
���u����Lq�){Z��Z�.hd�A���d��`�&�<$=9��wZ�������4��a�]�ޣ)�'-��8� �X��<�U����rY �&?أ�[��D
�Ie�ҩ��t#bY�ȶY�s��)��8r��,��r��1�p���vWiBd�sv [b�C���L�d�[լj�LHf����Opi�9��#�43V����n�vs�VR
K�����8�-��y�����w-��/ⷧǹ,���ޣt���X��lª��>-�5�f�(W��p��ACU%QM_��k�����d:}ߗ�e����� 6<�fF�HC�i{��1�s9�,Q!Ǜ�D�!6sb�"��3l�X�A�b�׬�
�h�����q'h&���TH-��Z�g���f�RH���d�"��Q�񛿓lsD$���A'5�֬ؐ�+Wx:�6�:K��[2Ԟ��G�лނ��l�����r�X�z�w�A�֦,u��h���P7�l����v�(�� I�k^PG'$����s�?�nY������z���pD�В˂A1`T�Z�����o�qy���[쎧lG����x������-�c{�>1_qA�}����ͻ8s�n;~/�N���'^�g&ǹ '4b��G�� �I� RH���1�k���ee�"�S�(��I��U:SIe�V���"��,f�6��:�Y�%W�#�nl�H1���(�_>��s��Ws�īxd�%�=�
N�|�%o�ũc/�̭/��ɗr��s8}��\غ�����R�S�	�-rw9( KA#2x��x>���<��|H��OJ>�is9W�Ƌ2MQ�H-�&�M�tzNg-�;�8B�1��Ai\I��E�ú^ֆ�j�7��>!eZ�0�b��p����H��!���ϼ���jI۔���5Ƶ*�g3T��
�c���>^AW|K�&��VG�Z�r�����;>t4�7����(�vťw���.�)����x '�`��_�9K�y�ˀ�$���`�q�����)|dԂ�V���v�����Ǜ���籧;�v��7�W�o{���g�K(�SZW��}����U 3�����9 %@ڿ��"ɏ
A&5^9��QQ��=��$;yƵ(8�u�<�GG�i�=��DP�%��02��p"��,S�f��"gO-5�x�r8�l��qp>*Z[�;8����\mri�ť��1�cA�o�M�yzǾ�<G�T�,��:'�s��h�E�#�$�5�����i��J��B�aS�����l1"eF&QIfγ�O�	W�On��L㹒8/
.�S.��c�eN..�cNUk�&炞rU�q��sdԌ�����A�ʡꨑ*Gg9]ptRbD`�#�TP(�	2��T�1	2������%W-�9,��,Y��>���>Ġ����
'l
�˒gB)��}]��*�/$H�!W���xgaq�Q־��1EE�v�{����_��tJg���
������Pw/%.�:�B�ÿ�&�����|)K<A�c���u�Dw���ב?��e�7����������|;���Ī�v��~	�\Q�w�iN���͑�����Y��im�9E�#�����m��-*4Hi�v�<���7����n����n/s���-G�vi$�k=S�P�/�#A"�!������a���<6�1�˜R� 6�]�� 4V���� �	*�h�!T�L&��D��(�����Zpvd˵|�kŐmYq�s\3����|V�(�Kj�Ǘ��.r��d�)�q:/xX�U��E�<OE�c�(ȵ�����-B �3�T�l��h���D�t�R}�Qᩛ�2��$VZ2��a���B%��*FY���|�8]�5�(��F������SΨ�sJq&ϹV���1WʊG��4��q���II�$�,� �X9lޡ�'w�<Jr$���̰*ê��*(�XY�Ba��*I�B�rE/���|r�b��^�9�m�yb�ِ-zt���qv����h��{�� ��C�/B��:��x��]�u��з=��	�i�y�1��Ǩ��
V�&!���3�j2�����`�U�N'�db�F��ػ��/���K�;��2����������tհ7^C�쵔�� 2�L��{�-NKp3��E&�E�u%�=/b�������O��h߲�Jl�F�c�֨��)�_��l��������x���#�J��>|�#��������{���h�����$�"��|_4$k�T�L��p"U�1b3I��,�:��Jpt%9Q+���-RI� (� ��4A	�(p���.�z���Ƅl�TE:�,X5�e�ɏ GG�����;�e6Pi*"��3	��YT��qIQ���]��|"J)$>���eY�dN�ζE�2*�X����e�S��4Z�T���0��ɼ@v-�EJU�:z��F�˖�Q)�� ��Z�SiY����2-���cjj�
ɤШРu�5R�	l�T
J���`hU����$9���L���O�j��G(B���$DgR����b�!"��:O��F#S���=���6����:a�KQHQB@��z.��Hɵ��@O�=r��_��ȃ�DaiT���;9����}/W�0eE�"u5`_�x1e�x��ۜh�Y���S�M?�'��/�4Ƿ�%�	�Ϝü��0���k#�]����4%�K�@AW	d&(.c~�L�%ˇt�&���?��3��C��g)��R�&(�/hl�w:֔r��]�O~�O~����o��d=[�0������>�Ɖ[yő2CZK�R�UAYh�G*(�^�X.���yO1(Raj�֥���L�[��bE��u�&�ђ�2�����u���4Ѳ򆦮�4I�F���s4�&`SЁ���ő�e�Ԃ=�E� Ɯr�QX�#��$��hM��й�؛���8��2�1ΦZ�6t��#�%G۶#��iZ��k&`lJ]4�цH':�r���[-qmM�c�t�b۲\Ή1���6|��ޖ�u�}D�1���:�R���f.=>E��	X9K�:��}K�Zd�(�l�Ce�LAN
N΁qd*Y�� ��]�8�Ip�n:b��E��ʂ�1�mM���,�D�"�� �4�.�]<,�������p�[h�����{�z;Y3Cdm���ο�����{�g�{�I�C�s(u�X�3{ds������W���]|M,RX{����˵��i��*cD*S�@�~����7ڮ8���P\ ���m��5�ݷ1>y�+�������%�ڏ���t�tk�l0F�����@��ܒ����w�8���|�����q���nƅ��&g��+�^���1��+F�Q8��`&!���`� ֑�xD��$�֎q�6�(��$W99AP:�*��R��:e�9��B+�*�1��u��,Ag�A�֒�.(rE�(Q�[��kjLh���am8f r�L1,$����pʤ2#ـ�0�Ԫ���`��G6���F��eQPV����(�yN�+��$�p��'��*K���9��%��b41MX��Q�%��b\���a5`m2fP(�lL������-�r�**�1y5$�*���"���j�xm�ޣ����2+��J�@��5te�*1
����ҊU;GO^��/մD9��[2ч�'�ĺT0{w�pR�T�u����>�GT����q���p�N�C@b�!j��
���-����i#	y���%���%/&[;�ܖĵM^��W�{�1~�߾���s�/]�[\eo�Q��z7�>�f>���Μ�����_�:lv�Zw�� z���Aڶer�V��u#i^��T/z	QKDW�(�'[n��{G�]F�&�[¹>�%���������,lVgY>�����~������O����e��]d�]�};�k����?Ϫ:�*:��S�޻x�G�H���s�=S��-.^{��T
L����2D��e�5J8f�[��缌߾����EfЍ������u�]C�I���`ȴ&X�����*d�n�#D�s��9F���A5@yO�vhQ�Ȩ�%��<�64x�J��f��h%Й"f�&.����>Dby�,3��8I*��5�uTk��\g88�����*T��+�s���X,��*r�m�TI�EƸU���d�ִ��Rm�ZB���G��n&�m��GEA�-��B�n,�(,/���E��1(�<1z�sd�s���l{�PHZ�	�J1n�N&��%�/�Y�/$��!MQR���\��q�ɗ�����O�����1�B�!ھ��De�^T��+/ȋ����9�������./��8�p���x�~s���񞉔��c�����]v�;C�ar��}/��W��;�b�p�����Ƀ?��x��о����2�3���b훿�X�[����f�썌?�.�qNմ�g��X��[��/����m�C�]Dw��kW8��r�.td�%߼���!w�v�rz����R�(/\���Y��/�~l@1�yPcɑvA7�q��G�"�mj�6�"������R�ve�Uca���;V�3���k�2�k;��JQ"*��"�8����<���o�H.$q���9Y^���vȊ��3��(�ґ�֓)�
!g��]��4�'c�V�ƃR� ���<�k�H2&�"'xO�u�Ѻ�-��D�{�"C�t�DTLgc�	6R�RK��d�CE	U�P"��%`�Z2VDA*LӠ2���"��.}�TEF�`��(#�( 8dG���¦�Z]�BGf}�'v�U�m::ћ�,�"c��6�Μ��+��V��QB�C X�-5yV��[���=�׶��cc��������7�S�e����k�j���%R��T�(+1���RIV�c�eh`w3�α{�eub���_���O�^�B�lB����#�ŜB�t]�1m6�[���~�7y�~~�;6A�[�9խ�4��P��־�ðD�����(#�4\|�;�]�T������~��\}���}�=�[�&8I]Li�Gy΋��<���5_��^�5<��ۈ���r�%C�?�6>�O~��o�M��ٱcL�����Ů S�c@�56Ը"PD�ւND���U�_c@����k�.�{�
�jE7_bVݬ��7t��`"M�P/�,�K\۰/[��Ő�n����$YF�yO�%�܂T�G+ɠ�R�s�Z�8�@H�/\m��{hdן�楡��9�[2�R:��D�:����[*bmGt�:��Ś�h�mQ:o�M�NS#`��e�$8�,$�v��Z����:��(]P��ΠBD�Ii)�'���m]�u+V�=�sH��ꚙmifܲ!��:v4X�n	�C���e�#���tx�\V{�=�s�΂����"����a�IG?z�7��q��!��{;���e�ɗ��r>���>�46��J�H*t^�4� �X�Ј �Υ�א�V�XfU
޷����Pd�QK}�О}�٩��z����G�?'8E5=����r��&�[I>�@D�H*�v�����|���>�+�lL��c�jI�$Ja��}%��_�$���?�� =�m���w���G�]��HpG��;����wbT�NG���W,�fn:tWCrS����$��%.���q���H�_�wC����J�F���Cf &8뱾�� ��X������&��ͩ2I,4~eh�t��jɸ��8/Q�#2b5 �DDDC�%ەCKX�c�O�Ȥd�����[��,��Yt�vN����c���t,�����س���}%�m3�a\��`ۖլIQCJ���l�&q�R+FUI9(����LQ��\�x�Zp�<On-S�\�$�ՂnѰ����J��a@ɨT���w�l$�AЬ�@�1���mBi|PH���AiZ
��dAd�\�BE�L�L��_V[��+�s�[��sg�]���.��9ށ��h"!��%�d�NPK^�4e5��X)�	Ck�uP�¯~-z��~?k�%��@:=-�!�L��z��8<�W �%�锁\eD,�Z�� k���d]�PA>��s��?�Ň?Ip-���|:!dd�2�$�r��k��6W�]~�W8�/�)�g�{"G$a}�|��\$c�(܉+j�{������6mBP�w��?z�>� YX�EG���xD�d��eXL`��_�}��7P~�W��:��RA��A�JB������������)v��1X[� �P�mD�i����.��u�T�jT�<�'�eP�_��o��_�8C���m�+�k�z�1�~�^��(�E�����u5Y���dP�|�k����5�7�LRf%^J�`L��&�3�'+22-��QJƣ	�|�|a�y��c��8�"�4Z(�sB������dX�r˭t6�w�,�ӵ��Ae���&�)����*����%�є���Do���:��g.20�\dm}J]7�F8�1�a�D�(Kbp4MM�	q�0�K�kX�,g5]�B����:Ad8���]TT�ȹg1�em2����<��p��GX-WD=fe3Z1B�&X���X	r[�b`z���s�J�1�/'ܧ2����=��u>��~��l�j��#W�qM�0U���b�
��$�l�����<g���i�a�3F�R�d��/h����*%�o�w���/���6�u���\��'���ؽK��ܦGģK�p9n]q��6ڋ����\U���'�؟�Q���.Z%�V�x�?�An��G(���j�f��nG^�L�
w�0��6�Z�-[��R���#�̡���p��?��q���C��ё�ǈa�j�����Xc��U��Q1ڈ4����>P�Y{!��9��k3Bu���K�]{�F��i#1D�"CFGN)V֒�r)H(��<�8��#G��׿����Ed*1j���N9s�
�r�#G6)�A�*Q%RB�j�s͉��9s��_����r�(�5�U�'�錦�t��)������F�1�{,�TÔBA+A�u���6�d���"H�1�S�:�T9eY1ߝ��1a8�Z�TU�q���t^!D�zO�4d*��l�1�#[�v�v�_>���m6�l�s���kj��<�m-�k)ˊ�@����iT4}Q2׵˒3�<ʻ��;�9}!ft6"d�5s)3�d�e�KF��d|�8[w�ü��VW�?�w��?�������lݍ)cK[�z��U�60�q+��i+�����:J���ɥ#�U:G�W�^`j�m���2�S�4�uj,5t;0Ca:d���i�%F�lqek��%�\�����+�o}G�؟J:������� �֜~�[��/�c�" W�4[컎��%㵊�$c�(Xs��G=r��m�yχ�N=��;?���)֖-��pt}������i�a�9env��:�@���T<Yi���Q�Y��6�!e�d� �!]����q.[Ů�L�ce��\�@<d�{�1�?:(�2�*5� ,*�Q����,��[q��^��X�ؾr��Wϲ�}k��̶w�5:�j���+'��b[��5�\�z����v��q��9�^��b��xT��]h��\�|����zm�rPRT�ѐ�p�h<a���eL�ʢ�9e^2�T#�dc<ec��ᘠ-B	Zۢ�*4�Y�(��"kk�kc����Q�������Ԅ.�>ݢ[Ο�����t���#�8q��2OR0(����x�ŝ%HM��u�zţ�α�#y5&�3$>����̩���rJ!�Ρ�$ �՘r�N������so�����K�}�{��B��2:��tYɨ��^`�F��B�,��e�7Z�|��
�$�R8���8�ba��<'��	�昀����c\�p��)ӣkl�~f(�]�͇�l�}F�c4r�sܴPLp�MK{߫���Pd��1��^]���7�����A	OX��{�L
fn�����%2�@�д�Pat12�Kc�Y:Z/J�u!%�α�E�
�US�Y%R�|y��+U�� �#c�AG"����Խ���+��&p����>�?��m��'��E��A6����iDL�8!�tF.s�<�e|�k��c'6�N*�-Ξ�{�ess')�1�Ւ�y1 ��֒�9!F>����c0��6e��Zkb����L�����hB6V�`�:��!$�ф<Zj:��O5}�(���@���1v>8@&��H���Z�Ne �x�D}�u����,���Zj�RH%�����NQJ��kB���3���Vu2�e�<�R�u� �bt����KWNs��6o{�ﲻ�0M�ݒ�����.��JS�%~���-��7����wіc��9�����+����vν�_p��5�dܘ"�Yb�&@�`�����T�20�迸1`��o����<�D�Y5+���S��CT�
���2���*��Fe���v�c�c=*���l�#9�f�&�3�M��d���S�u|��숁�~+�����ƈ��1�=�ƃ���<�`:a�u�;3v�Wɋ]�D��YVaf���б`oU�,4DL�����d̢��P��e��t�U���6���Z�! �$K%�H�	>��V�d��\��ͧ�|o�w���t����;�80�d$S�T�#A6H���0VR�����K���k���/asc��A�bY��!�`H��Ūf�X���[T�!�GtQ"��� �5JI��!��@bRZk�4MJ΋�?Σ��1 PZ��DE�u見�&4 @I��k��ާc��e��\ؘ�P�a���pE*Nޥ*o>x�%�px�Rb��޿B ˓�'8C�e(�p�b�!���%q�]@"�6H�z�
���C��/�*;Wk��:�G�PS�%����!�JiB�ĬT"b|d��	N�}'��eg�U��?��<�� ���|���9'D���h_#�N���ꏒ�2�&�;�5�� �xkQ�!%�3��&q݊</i}���dB�Z�ҙ���_1���sdYI�m�(��K�|�Z���$c�b(Z;����y�x������W��&C�����Ԝ{��)���XP_ާL���ML3�Cal�tr�zoI��7�i�B�k���HTQ���Xg֩�*Ŏ*M�;��,f(�c�A"���f���іngy'���K+����N��9(E����ƍ�6��6�`�l˩������p�p�1��1ȀdPD��H:9�Su*��+y��Ƿ�1�ء�X�֪o~s���<��T���"�ƸZ�wW���R8
������'�
��Ѳ1�:S+O�@ؒ��$�Gz�:�%q�x��y��GYZY���c��H��Օu������X^��4��IHZ1I�M�ĭ���`ا?�nw鴻�0 #�$!#� �����uI�@i"�D	Zi�(!P!�T��Q(�4A�J4����Y�RG1I��UH+�B ()	t��� %$Q6ϭ�vBj�R��MH��G��(���#b��-q��q���sZ�D!I��c^8%	���K���Hd#6w^�	�5��@Ԙ�DX���,HIk�a��LI�7�X(��^���w�`����[*A	�uv�&Ŋ�Am��ƅ��YF�$�����֐G-
ƨ�Kjj���QBja���)����b�9��!���t�'���6�Ŝ�,7Cī$Y���ܺ���S�����}��5�����P#��X�@y20�*:�'�K-���;k��-��g8y�zĭ-v�d-�,)ط
�`G,t�	c
c�&8hM�R�/�`�z��,!�=�� k=����}*�DZ�9��)ʪM�AeZ�E�*T�֥��uE�R�ԥ�ۚH
zڳé��l�qN���#Θ=�Ò�,YN$��sl��0����V��p�$nF�v�n6�O�x�� l���#əCE@�B�ɐHF�8C5_+��B{Gj"-iE!�V�"-	EMx��jC;Դ�&���Ҵ���5]�骀D(��ha�!RMM�͏��5� �m��ha��o~�tDʑ�H@ ��XI�քJ�q"�G�F*'�ř_�4��3�PDk+˜Zp�㹣�q!8�8�SM�Q��m̢�4]S�h T�!�u(�4�@�X��`gg�1 P�c����ZKΡ|F��=dw��P1�4u-�\H�|�ò�0P̖79��px���)��'ُ��),zg؏�XtN2��12U �,(���'�mA�d,X`DI�Tw^�<�ʪ\e6��	�3���Ü��f\;����5�*�G����JҚ��?�<p{�v����撘ӏ���)���-tR9�h����� 촑��$h!���DH�bF+j�sZ�B���ޠ��bJ-�v���X^�Si1����h<��}!�`������KӔ,i�$��w^{ku�F8E,q�qlYqv9��a'8�`�� ?�mLr߻>��G�xA�j5Nc1�����+0�k�B��-��EkMō�D$��(n���caԼv���H`�	Z=��CD��5z�uEJ���7� �UE]�(-�U�s� R'mTam����
�i�3��X'�:@+����h�L�," �B�#��(!��,:�Q:$+*LU5G]�ȳ���z�5���0ƠdI��9(�S��.��ȽWiyW�f��q#���aHA�la���6��-6N���Y�Hɿ��������yB�y��l���(YceN�deg��n̥��]�'���`k&�f����T5����Ǖ٘@iB��9R���ҎC���
A�,e �֎~^�j������Y,���R����u�ԯ����߸��,<6�P�֠?��?�S���C�Ϯs�Ȼ�����cD�-��d4��Y��1��\�S���������������3硶��_�itD�I+G)Ӧ��4H,�ToQJQ�t�4���$���hE���~�?�?��ע*.�s�s�{7�a�Q�-�~�wya�E�:������mi���Uʩ�;6ڴ�.�����d�W�W�q��ztw�钕%*�u��MT�o=J7u�w������()B5���7y/�7�>!�7�^-��T<��E�V��M��g��Ci�(d=#��k�@���%�v���*UU��k�"E���yIm%U큀�j$v�FfQI��H���?�Dc�)��׍A��ZK�֔y�������ZP77Bb�Y�{$����6f4��G���,K��'�$�yM�1��`�'��@�b�r����?�W�3|�F����_s�b�	7��S�$g�Q�=��P9��������W�}��.���i�0���~�Y� ��6��8��(���c��X+f*Ɩ��I��x�  C��U:g�x�c�����_��`Q��	z���_���W��q���6�=������������'>�I�@9��~
���\����E���W?�������Q6z�g/]����0s�C���!�N����dĮq�v��
�U!�xn;ɶ�y�c?��y�פ���f�̊��Y�[W�S*ŷ^~�K�{���[��W��[���lg�7&�Ld���	�+���(HG3�c�E*��5�n�`��K�j�w�p�<r�,Qo	:��˄�V��'�*fy�5�E=�e��iIZTd����S+���E���BRV�� D��%i)��N��E�	(K�U`k����4�EM:�8�Q卝�TH�;H�È��5�hn�~���I���YZ3�̘/R��R������U�w
)#���=���2B�	a�!JzT^��X�uޅT�l��2$��#�IBQ5*.kE3����(k��1u晦�B&L�.�O��T���N�$�����J�S�^�^�G	����^�w=�o�q�È��=ͺq�*���&(���ß�;,����4��l���A�������cQ��+���h�գH�N��"_���RxR�n��$$�D����faKJ_��������#���w�����*9=X���\y�&�����7��hBt�C����_��'
]�����ؙ��;��O��٧���U�ɿ����a�{X��"�~���������%�ٹ�HH�Ǡjѭ��m�h{I���(��9Vd��	h-*�j���X�%� &�:�H����������=��<�����l�y���x�m�r�T�ORr�|�p��hw;�VW��!��E>8Ǹw�K�8�a�9�Cf�ʹФFc	1> �\���P��T�;���P))��HE���^�>�r�J�p"$/.��2����W��ao{J�Daİ;�7Xfi�D�7�'�Nr���l?��t8d��y��1��qV�NciS��a�A�U)9<̙L-U�����6@�S� �5F[J	��)�#u9��\9��Q-#��D�PABa<�
��ܣqh*�V����?s�d�!1��hq�ZTuD�d��L��(�=\&��Q�1�-Nz:݈A? ;""R1�}׻�ꗟ�w��3�F�)e'������8���[�_2<�|�������˅�~��Q�bf������s���3�(�K��d��1ݕ�EEET�gym��(>�@B`$}3M�#���������}��������s/��N�#�����ϣ}̅S,=p"�5�kRL���x��9�(ldX�czAëO\}�Y>��_�K���|�WXJ�	�bZnȁTL�	Y+ �$VK����!ZS
F��0��̄���CAZ��8aD��|
'�y�/�8��_���	�8��x]2��}L���|(�o�	�H C��%Q�&�[8��kɭ��f*0�)��D�!�����ؾ���b��>�Ǘ{�zD�أ.g�ł�N�֔�!.c�1�)���:E+C�N#��q��k
4�-S�s�NA�TfNa3�E���R����C���8q��`�g���O~��w�}'����w}����&57w2��?����]<������#����<���I�%�{+�=u��gϳ��L�A$����Hq�{�����yI1��*UAhj��eE��A:�:�2)^T�����@.��Tx1ao:';A�Nkʍ�y~��|���>�eEmr.�E^�f2�ÙA�Y{b�/m-p�ŔSL���%Zݚ徧�Y�ᰧ�fł���EHKo��C����.ɱcxb>�_������ޯ�!	���ϲwk�S"ե�#�0�*J�}�"����G]�ĦDNXL���Q>�6=�$#��u�z�:;��Ez8e�F
�T�����6rWQ������!���?�I�&�=�W_�p&���Y�}�9��Ұ��;a�xo�O�گp�޻���������b��BQd(Y���z"%Q^4]Bg�F�&�D�%ԎDkb��x��
n߼��_}������7�Wx��9�I0�_ �z�������0�k�9�h<��jB%�}��"��A�x�g.%�����і���Ha�����8G4�{�F��"��9��U]�Ú�.^W%�m敦i'6V/c��a�f�h�&�4C�,�Y��f(���X�	�k,{���޺|��{�/~��y���O�e�˯�ɷ�}�+�.��˯��K��ƛoq��m����˚0�W�0hjPS3�s��D���nLcY���|��U���b����TXۼֲ2[74{�p�P��xW�1D��6��.�� �Gx���Ǭ,���Y��Xa��iKEA9��*K$%��e:�!�Pҩk��p��~������9.�jS���'�-�C��yb�o������ν�C�j����?�ﺌv�,�f��7v��:�H����Qx8�tR�DJ[I%&��l��#��J������)�1�~̛_�Q7!ZY���x����/s��<p��/1��?��#���;6B�.��!󘝷)��t�q�y�rx8��;o�nw������ ��Mf� �EN�Xڕ%tY�hS)�P�M�[��u��*DiQ�#������?�g�c����q�[/�7�n-��<7f'�M���Pň�:h�� *�AA��US�-J�t���.;儉4d� s4Q�������XLY2��HӔ��I��<�n��|�4���ߧ��u�Gv��|�|�`:_0�g��f�)�,e4����̦s�Ɠ)�q�Q�=�Ɍ7o��K���g_�_�p�aJ�d:'�Μ?χ>�N�8E�Nx����E��s�W_�/�)v��.c�\�z���|���{L�3��)�b�l:c4qx�<F�1�ɜ�b�b�`4���9�iF�eL�f�9y^㜥.-y���͙�d���(Y,2�Ґ�%Y��������:�{��S7�߭ �t%�lFe�RU%�Tĥ�m-�,��T՜��UL��W���My�u���rp�`|8ez�2��A_�z�wH���>�����]����,Q[ǳ��c�-�B�����!��HA'	�RHz�>��-�h�
Zdu���u�:ņq_��ڏ�#?��h�SOޠ�� D'��Z@�Q�!��n#�����~��QZ��g>�;��;Or�k�O��5x���w)��y�m��;>�ko^�o�N'�#�@#58��@h�<���4x-�J u�\�P2�(�X|Oc�ᎋw��7��*s��!d9�Ă���:͙/r��͍���Ī��DD:�#�CZE��5,���ҵ�D��I�_V�YI8-���iV`��Q�A��X����
F��d���3�<'/�<��J�2�#H��<ͩlE�VX�ʲ�E���(H�9Y^P���<����;*Saj�d� �*Z�.�k�q��|��y^�ڬ������}�y�2�x|�a����?��������i�x�qs{��|�t�c��2���(���b�b1g���u�(���;OY�U���9���yOY�E�"KI�)yQRV9�EN��E�l2��s�,e1���E^P�Ŕy���f�eY�g�*c����e�#�
��N�!����1�E�œ�v5�Jp��W����^J𵠻���N������Ƕ�?�k/�և?į��5�w.3�Ա' �>L��Evz�QŤu����8�p�&S��4$�V.��/5�\Q3����2�<��O�SW!>�X]:�!����p�ʌ���o>�5��3�>� �!R����v�{)��i!���8}�+�]Z��Ҥl��~���[��RΨՂI�M)��P��5�YCB�k�$E�ib��T��eȲ��f5�ޔ��,�+�0���{iN����'ܿM0�0�
�ft���*���ƣ�
�^*�T8��%�=�Gy��(f�iQS�9^)�N�N����l�����i��Um���� J:̊�	a�Q��BDQ1a�W(%QaH�B��}�v��
���*���eYp0��������·�}��޹ƕ�7����\#/-7��y����;�۟�,���Ԅ��ss{�9���c�Y�<�SV9I���:���n��FjM��I�%A�N:�6:��u#�R�8nH��"��Sde� bP��8
��n����mҶ��4�	*kȜ#��Zx�#�Zy��}�o�ͩ5�O�yx9�a[��bFRUTׯ�hD��.[dem��h�;�X\�a����K��W�EG\��E�(
�ʠ3K~�|w�0��r��~ʤS0�SR*�0��0�K��G�1���/�������h��|���b<��L�],��I�L��T��ٿ�I#%a1����7rm����z�u����,&l�y7�	U���7�ɫ����>G����P����.�BEU�~�m�-��ȨA����	��|<��+�1��Y^Z�:Ϣ�)u�;B��|��`\��؛PG-Tb�#�N0���X'(+K-%3<�@b{]l�E���Rː��v��V���<%��Da@�n�kJ��t�T�4R(�H��;	���A�3��}�&0E
oJ��x %Bzz��3�(lHBb�!�+��h���xĵ7�ǤY�����|���7n�Εk���������R��+7n0��t{=���g�$�EqL��Fk����jrG�'P�<���x�SW)P*hn.A>�Q�D�p�Q��͢n�;*@�$�	�y�ڵVH�� N�8�A�	ct�)���L�]_#�t��Sz;u��`2�9����W>G��s"P]�AǄ[����/sv���[L���G�q0��{��l�Q����õA'�+��6��xW�us"(<*�����p^4��
�a�ace��_���D�Ex��w݅5�\�x�k\Zx�x������$��l>�>�����6Sc4!:T����t�ýw?H��B+p��m������:�\B�>I��t�i����P�@[E5�0iE[&D*&�b�a���k�\:,M-'kϠ?��Lgs� �%A��Z[pܿ�-s��EejBJ��P�ysYM�Z�Qs;P��#�(���E[��MA����v�$"��:-��>Z5zRS;�R�:1�Kt��B�R*S�@:�s�:�9(f��k�u�D� Cz�� ��wc8J�jutТ���7n��X/�2��P���w�t�
�yF�c�����:E��:}�iI)	^�E)����(u�P�(M\`qX_Sy�V�0NP2@H��b�H��8A��TGBI��a�0|���r�p��W*����#c��("k%LXOZ�m*�s����`����[;����p�e��
���W���Rj���̱;�Jβ~ϣ���qz\�=<B%���2u9e������&Eɼ����U[b'�zE�����n����4w�;K��͒�Բ�,�y
A�_���O��?ʕ d�M���Đ�{��*�,��"��{/a+�~�Y��"����:w<���\��3.�6U���G���v`lN-ԑ�j�Z@���s2L�jC�X��ĝ�		ֺS6�:�C}�?����ǐ](;17҂)��fT�!�GKA [�i�蠋��	dD�)z)lԚ�j"B���l���c�E8��d�襥�����Zĺ�#���]4FFM�T!q�M��i���/E�'�!	8�A��QZ�T�8T�C#� j��Pk��](�Z�Zm�v���A�Q$�ۥM��CF�	IM�<PR�P͂�B6]F!�>D:�W�"@j�
��-�ƙ��;�VQҢ��҉;��m�R͉I���^	�T�@��jN��>�X*A"�&�	��t7�h���)C*4��c5/898F�L��6��?`�K��sP���K������7�]�>�0�k<�����_x�'�+�<�"H�5��cܕ�؝�۷�ܸ���kLw��w�u��%YY1]d,�ˬ�����;�� @꿂ۇ��8�a��e�>|�U�`��a{��挞�P���A;j��G��������:���~���������g�a�����_�2���uX^&ܻ�R]p���W�±0���j�Ma��Q�������/���q��S겠����EF=[в�NYsgo��Q��ZC>t�N���|��*o��>�q���v05�@H��)T����X(IH�0D*I��#�b�xj%r�h4�J�&�45J��1q`���h.t)��x)�$G��5��RaqL��F'R	�lw��ä�pYRXٸ��SR��ȉ;
�ib�H�X�����Æ�F1�8F� %C-H�i��%�K����U�\Z��Mt��Pj�nj�(�� G;��}t��Z�lH��[��8G�������[�e.<�I8�|#��YJYT�Z1a�mu�[1���V9��?Ev�*>�9qz��S����ͳ���:`P��Y�������o�������y���S���3/ ^��t{���ܞa&3�8EL2�lF��P�j<F�Ǩ�5�b�#�tBr8&�?�O1{��M��5.$��u�)�xO���|�S����5&��Ϥ=��w�˥�������q�{�D�����R[��&�<���}N~�����\z�e��������y��_���"߻E���d���]�12d��COI�h�����9z6C�f�ل`1GN&���.6/���"����fU*�7�Q�ڥ���~4q�`�Ea(�&Q��yf�)�bA���
���U��!i�	�-2[Q�TE(�Q��RM�$\s�JD�i����ԑ8\-�0���M,�sXg�4M/܈�ASwI�y'�� Ѵ�]Za�9�G�i"i�`��wxDs�h>���.E����E	�&�N%T�82T�DHE����G�wq�q�	J�&`I+�DI��=���'��b8_�]3ӕA��t�$8�3�*����M,_�,ms��"����jaʚv� CM!��r��:�;�н>[w���u�
6�V�1��Q����iՖ���d���w0ctU0zt�.Rh�4x�(�D��@Jz���zeŒ���vZW9�)Ns�H������6V�8���iӉzl��9~\S5<x�����;w����-��:ϱ���"[�>05zv�������ߛ��;\����	�wn�[^gx�ۯ]b��[� ��^��h�r��uF���r�[W���=`qu�~���%����U	6��CR%0��vq@�R����뀡.�-m2r!g>������
_�拈h���͡��y�6~o�<���S��r��L];fYA��1��5�bAM)�2@@m��.(��
����kz��\�j~N)�o@_:p���usaDG����K)��uM��yN����3T�
=������<H���I�h�i"~��G��v;�*�de�ރ@"����HJ����G���{\]�f'�	��-P��@WZa=8��#d��cLcbj���j��5Nz��H-��Q�)A*	F`�EI[�J(di(�g$Np~��ќ�3�P�]nUs��_x�y��x��{������O0�w�Pަ{k�����ϒ��V�*g.|k�/�Ӕ2�d�xo�Q6k��;������y���%$��0y�m�_��.y��g=e�X5�ܢￇ��>�A����N��]�y��a���aU�2�*�#����V
��,���y���o(�1��� �����;3;�3���n����/���⒐��_�Ǩ������9����~��@k�]��_�W����K�@Ovw����ۼs�:�Nq�K�i4����\�Р���,���J�L��c���KB���u�(j�����K���{{Wy��6�o7)Q�sp��[���.�4'Br��)�xJ��Nz�s#���;��7�@ZO�Jx�gP�I���BЊ[��j:��`�G�[9��8��&�v����߻?z^�ԁ�G���2�A+���<�(ƀ��D� ɛ�RJ6GS'�J�Q8_#Ds�7x|�+��8�����G4���XFԮ<r�4�(�u�|`]�[6�s`,����		r�A�O]���&@�&��4��<onr2)Xq�R{��5��8�s��&�Ɛ��::J�/�[?����~��;�������qO5'	�2C�t�%d2��CP��u$s'�U�c�;��O-[8�aZ��{�:�,�^s�Gy���(�m"�C
���	k�
N?qO�z��t���	���%@��*v�:��=b�Pפ+k���w���8}�*����yy�яq�_�	|���ә�ɐxt�w~�_����c�*HN�����7��0^fQH�����g~�XH���9�rx��ʸ�el���.]�ItB�Us���0���Aw��1�Mi�!�[B%�@]ۦ�2Vâ��Lֹvf�+²�T��0%7�_c���q�v�H֥b��TYF�����S�"��4�F�D�^ �G�6!��8��6d��V�qP��s��ت��h��<I+�2�'��� h�2B7�>�ZzjS�(��ޠD�W�GȒ@��MX��y4���D�څh��VZ��x�V
�"�
�w���p

�����W��!d�mnR��U�����m#El�i����9�P�}��Ch�w
%�6�q'$^X��,�j	���T�I�w��3�%ǖX����K;SN'����!{�itg�G�sO}��x��V{G.*BQO���dZb��(�Kd��	�ꂎ�-R4�8�ٛ�1�%���O�v�Bx�P́ +h/:kmD[SI����E YAt�&�����o0x��r��#�=�~�����|���O<zϣ\�:g��r�_���~�?��O*׎+_�"��[�'d��D��ͷ9#"�!���Y�KG'��R�����X:�'��9�:M�Y�y���k�N�Ll�x���8�XE�*kb'iKE\V��d�IeY	5=�Y���k�!��gя-r�
D(P�f��5�r%э#��_dRh4�S�$@Y	�"���:��M���@"�o\�Q��ġ"�k<q�� MS�B���'dL���G�h�Y-�5QJ��<�&�Tʦ��&P%4R�F��,����!�.��]8��$l���fު�@!Ax�h<��5Y*B7�h֝��u-�	��6��#�S�U3f	�S/���L܁�Gn!�h�+������Ҡ!)-�dFGV���c�Α�5�IA��s�7^}�LG���E^���U�4K9XdL�b6e��q�3M3���y�h��0�3�k&ل��S3��Y�)����)��Lf�3<}iI��]o��j��vhg%�Y���'�^���k̷o1�kV|L8SD�\9f��)��,br���Ӹ����yV}�����JǴ.��Jn�+��!�>$<S9��^A�cr�\�V=�*���/1]L8�u�0��6�-�� �AJKLHO��ɀ|�Ŏ�����L'��!�nQ����́vL��lA�Wă��ed_��9O(8�χ���U��4���@hZa�A�pE��BiM�Ry�lR��o�3��p��T͢�4��6/�+K�#�P(�o:�h�>
S�B�ćV�E�%���]"��4�"�4&�HɆ/���B���-����2"P�H4pd�-x��U��DA���i� ��[5��#���[	O�V∅��A�4�UG
Tp�C��|�����t�+s|]�ŗ�P[��B��ê45-5�xdm�1ZJ�A@�5U^��g�FX��x4`��C���t�7/�+W�xc^���7�kp��|���f|�J�KW+.]\�%����rk�Ko����W���r�6������]����H�}�`�G��(n��{�
Q>A%�zɑs��p���J8�L�L@'�C��k���yXT�vR5� !P?����I�*��ųϰu{̫�B�y�;�]�Q�7xG�,=��!A�bF�/�~����a�+8:|��7�z�=D[ǹ<��6��H���B���
�W��=ZC�a�v�ɦ`3��W����Ȋ���щ���rs4�0��x6�0�Ψ�G!�CKI��S%"�Ȗ���m�-����H���h���A�a���P��4
(i"��X!�V@�t0�T�@��<J�4B+�VR�������2D�:<:*��^�4�6G|)\��L�
�Z#��X������I�r�C�u{�*E*��a�!�0�5��R�����&9��ϵ�뛨v���DD{!P(���̊˪&n%B5��#�����o*y]��**�t�fw@7��.���fSҲ&��;ϱ�ⷨ�Vy�C����>ǉ~���q�>a{��֏Q,����on0?�E��I�qs����� �~�ri�ŠO��
�ϲXY�\�`�p�yn	�����2d'��9\��`��,-�V�W�C�&<o�7�?���>��AYŸ��nk��w��r{VrX�����Q�����#� �1)�2���6/��M�3Os��
�O����)Ci�9sXל}�>�K�0��ǷZ��j�7Op嵷XU�K圍s��9W�\'L,R�ifZ���F��%Ȁ�9և=�)�q(�j�I;��h��y�8I�2A��G!��]aogJ�0��N�9��ev�,awH���c=��s��_֛�j�@��r��	�UH�	�����`15�@�D!�<%J�Ԧ�[��� �kH�c��cQ����kMs\��&��Z�Զ�U��(�|�U��Usc �n�C����^�[0):RX+Qʣ��x��ڦ��ٯrMCH��u��NQaP�7�<�8�u��/����J5ia�	�5֠d����:4���P��`<C^�宍�I�5d徻�2�q���N�����n���O����ڏ|?��7~��E�O!em���w fk��}�CtΟ� K�|�x4'Jb�2�$��[7x덷)�k ����̈���I��4OQ�E;i1ͦ�{�'S2ȅ!*K��7�?����;��,�q��w��S%
Ο��o����&{��{��;�����_�N���O��'�U�(�|�̛�Ļ�w��?�tm�?��O|�Qҥ}�ڏ�����d��w��=��,���ig�'3^�K�`�^�0Nb�I�A;�VGs�%�օ��Aw�����v��8�Z^�|����{��|��{�c�]����>���}7�O<�[�1o�q�-zH'���,���� �
�4ǫ��bU@eJ*ie���DI�����n�!H���LSIj�xE�0�
D�����b�D�t3���lsQ�@��:��H�����(u4�ẀV5��
�GO5�/R5z_�P�q�$Dx�,4��TX�+PM�ԫB݀��F�qMMi��[K� �����w�]�p�a��I�zJo0e��4�]�)��{�t���)ф��f�BЌ�����]u��u�tA0����H��:��x���Mvn퐑�=�~7W��u���x���<����	���v"ƐT����X����?�w�_z������_}�7�9o�ؼ�w�{�k2��
yw�]��%C�V���f�xU�D(�2�@���Y�&u������K��LUwy�'X�3w>����̆�_�K?�?�*���?Ǜ���Ŕ��]�?�X�2������dK|U����.�D?|�{��O��o�
���?�ťK��}�_���`���3���sf�9b���E�nբgcD"���PDh�	rGPxzD�
K�.�T�Xgsbk���+��·���k���7���%^��Wx�O���/��tY�,s��5DtG_�h�(�Պ&q�1�%bsD��t�_B� �o*��h))�W�-Zx�tA��C���M]�$�5�DU{�vc	���y��h�P� "�\SG�2B	�0�CZ���@8B4���$$G��V�P	�whئ&��W͌2�L�R!���h@��@)!���SoIz���$h�N��P��P4���yB�VDH�@�H�V�H����P�!&y	�TH�w$I��WWx v�X
�E�t~|�D��H�=��a��s0e5�|pe�΋��;�Ņ���|�G)8�
.����9����9����,����o�}������7ޠX8k������.�؟pj}[Y�o�	I��i��j��}�xn�C�g��C�����UE4��H�,�1�W�����=���s��,�����w�x�9�U����$W������E�{�Y���;�����4��S_E-�x��$������Wx�O���?̅�>���.�=�ƃ���)y���&�%��!C��Ac�RM�"�A{���Hh����3��:�YPJI���][��}�p⎋�Џ����>�bow���;l�yZp��m����+���Q6"(=Iң���V��+����ro@hjboh��X4m� GWK�QH�%�*	�D4�XQWhk.�whg�����y�����4Q���B{����;D]�Y�`,5���� M�rY���FVE��P�)y�tQ���BU%���.�E�/s���� M�vijD�CQ�
_U���&�"��3l���sɪ�����Y�/JL���Q�Ȫ�����$u#"�Ƣ|�QW5�:��D�F�dk��(cH��Gt������X�������ڨHc�@zܞN���O��;���s��؇vC��_�#6�(�S�������i�%o�ҿ���䎏|��?�|�>�#�{�s�7�-���%7vp�@!�� �0��E5G �$�t�[��'��@��|^�"!��8�Ȭ�ܝg����9&�������S�*�y��z��_���'?�ᷞ��Vw����A�Q�����I'<z:��/}	s���>����+6W�t��w�=u��6X��bė���|�Wx��>�0$�u)�$j��P5�)�U��G�����--��Lj����M��鷙LF\�v��bN�i��g���ӝ]�ۻ\|'��ƛ����2�Z��f��a!0���n�KGz�E
����PX:ΣLE�P�P�[��A��|�+ң���d)���ĕ�(pY��3\�c�9&�(s|�S-f�iJ5�Q.��<�\��"�.
l�AYc�9u��,�yZf����qe�/3|]!�_U�"�e%�̱ق*�e�I��"�u�+J|Q�m��j\U!L��rl�a��/�)u�6��l�Wd��S��s_d�Y��s�|�I3l�c��*+����S�+�ܔ�E���C�&�WZ��+B'���8�ך�&��I&%�,i��H#�}���:����go_��|/�|�l��,E}Y� ��no�q�]�΋ϲ����"�d����΃������_��<��s,��&H$Y��P�BP�� �h�� �R�%jkQ~�&.��	�w$�L�N��x�ԏ�0������c'Є�[����iq��q닿ǒT,Μa��f�FW�"��DHފJX8N%�h;�u!Y橉��_���I<�T��6Y���[����ȒP��� c%�i�� �I�I��חa1嘯�����t[Pܾ����]ǷX�D���"W^�o~���9u��ﾓ�Ӎ#6W�Y�$D]�RHtKD!Bh*YY!MԼk��~�����)b:%,kzGE���QE���(MT�|Nd�Y���i���~`H�PI:ғHA�ڕ�o-K� EO@"*V:	����0l%�XZ�ذ����R��c��QıV�j+d)�t��/jR��h��1+�k툕V�jr���Ԡ�rK�E�6��ȉꌎ���_�؊�ִ�e!X�!=�i��.�e+J2TC-�KI��%-�8O��B�"<�R2P��@�J�8���mK�2GetV���������*[�3%��dYB�	�'�$�|AY�B���qrm��h6Z�~5"پ����x�c\8y�S��Ed%�'OaG���'>����U�`���X����!���_��=�t���7��쫸�B9I[�(���ܲuH\H(B�ܒ9�Tm̼&n������p|i�OG����K+|�O�ǭ�v��<!��`�G�e����ID���]N#��LT�ϸ{z��F��-�o�px�M��#ly�SC68�������>p/��*a7eΙХj�!�d��L	�%ף#�tRCk�q�r���Z";�(�t�΀�;`��i޸zZ}|my{/c�� 3�)��6�zH�!X܉V1���FLT�B�onRсp�$@�0���_�!%.���8K�DԢ��͔����n�.bd�}@�A�q�Z�!�8�!�d.pVᓀ"0̃�JL��eT��3Ŝ\��g{��)�5T��:��P�B���hN��66q���<cW:a@��(Q�#FdR��9)���%�%�^@ٳ�]� �!:�0i�-<�!8�
Ұ��}��ڒE�(0���PPG�#�$�JbT����	U@�h2��k�l�P�
J�)�G $��e��2�%\u%cS3+|�O��i*աĲy|��z��-ρ��f{(�q�f.���ls�5��]�nM�-ÿ�W�U��CkV��3_��`���̯N(�+����"l���Q,�eJQ�t�{f�dI�����1�+D�}S��Uo΋�	�I���LoZ�x���:�A9!*�,���BX�V"��
����2����$:���"Vy�7�JQey��
��<�L�3Z�^f�FO����(o��b0���S�Q�XK��HY��#���|�`6���L�� �9�s���֫U���6��U�������*���YX4[A�@E$^ъ%��ı#t؛�se{�k���ޟ0�+�$I�(�5Tu�S`�d\��t�F��*eZ�L���-��%���b)�G�C՞�T,���5�(�B�p�$U�E6g��S�|ZQ�M�pܢ��E�qRC��8�N+��GclU1����9EUSG�%�(�:�B�T3Fa@Ћ!j���X��:���7IY!
_U�V��<�1��I����������Q���1�7w�٭Fҳ�EUQ9�vh籵�hG��w��������/��ko]bgw�ʀl��]��F{\~�n��:��^#����`y���yh� \!�.`6î�����Y0��۰(y��יL����.I[3%�'�޲?=��Rt+�(A��D�;$���ۈ"#�5�-�/TU��+����j��.��}p�?��?�ӟ�G{�ٔ��C��y;3u�f��Yde�l��F�X�����Y�A�	� ��*����G�Uԩ�s��<o�y��@-
���9�:%1Z�(�
�FY��T�ƕ�*%kB�\��Ԙ4%=���nS�GyA�J&�=���DŌ�q����$�q�'��Jҥ�,���[�EMO+ph_�ME�-O��7vG\����hNe<���NxK�*rU��5����y�9hin���wn�֍�u�*o߸΍Řk�!U��V8�.�-��d��
A���ԝ��H�ғ(I�$2A�����!�Y��9�t�C0\[c8\��#ʬQ���,1�S���U5]��I����sd�FG!��5��1J�D+C:k�t��V(�)\M�,Rj�q��K��P^#t@^FY��x���}.O���8��t�a�R��"q�jc��fb�F��%� ln�Q� E�:��<���q�����u�˕�乻0����1y�2�]�tp#CK��!��1~�sO����?�Z;��`�-x�Q67����x�,��3��HV��.�q�d�+d+a^&Y�x<c:Z0�OQӌ��QuEUͰV�
*ř�����CV���>�/���7��=�^������>�x?���K���[K��8a�
*jgd��5�z�7�f����>`|y�o���_�o��cU{���%�n@�ה��i�;T2�H#	a�J�8��B�� [�X�wc��Ͼʭ�����e�;�<�{��|�.�)�oѺ�M�k��>���V�A7"5Jy���6G�Y���w�x���kl�=�/�y�a�%�j 4��(�\.8�y��x	�V��C���p���q7\����'虨� z�u �h��B6��8�V	Fj�-�]	Z"�tN���fŜ̔LmEz8!P-\�E�iS�4��(�&t*��� ���6*jS{H�Ņ��;GK5�.�&+-Ӄ�NHʺnНy��bJH��uElKu�?H�˄�'9�[��`������3wqgw��N�N7!
E�c�I�EQ�U#�X�X��ٳ�<w���qvu��vD(�
�<���chg��9g��k���9��,/��$8w���P�}�J��jL|�g�W~����^����G�}:��%]kQ&���7y������*�D6�K�YXp��L�mM���f&Ed�� 	4CS��3W`�)�#��d�~g���gH�e'��`�:m�	�ʠ��D�o+�L���-�,fE�`��6[������P3<���>�+�<��b�G{-!m�\�{T���O�T6!uVDTDT2����\Rᩄ&���jO�$yl1��{f����bεlFtl�{N����w��7^f�9,KLY�Fc�����7Xj�l�.��I�-T���+Oa�D��%+�ܱr��~��0f)�pr[`���_�TEEQ��Zsco�Y5GYHʊ�T���P�5�4SfjQ�JO�e��QbeEl���&FѱWd��CIkr-�]��e�$���]�)K�����1-
eCl�1vQ�-�H��Iੁ`VW�,u^V�
4R���Bb�a�,�Ȓ��v�E�"�CY�'Kf�e�����<��KRZ�GT�q�1�5�U��l�0L6�RS&
BOGy��a������
��Q���Ď���	F�~�ӧN�����|�}�Lh׆ ����X���/�6X���	�7���`aX^�`�b�~�q����gߠ>u[����?�h鐕�M�@[CGB[	Z��Q9�A�ޤgz�˄�hS�Y幽�ϸ*�1��������x�����0X[csm��'�2�T	2�����, �t�	�!�.�4)K�����x��	�{�H���m._z��'W�����\�WT�b��
tY�-G��gҕx��R��IlNh�DuM\ר�"�+�ib�V�7�<����
O<�.N�u'�y�7���=�m��P\~�u_z�d��d���ْ���e��=��(�(]�(@�1��t�dus���
�*��/��9� z�.��6��>B eH'�p��)�7�Ytѵ%@�������ur�Hgi'q+au�ݍ��6�Jc�AXCF�$�^���-�yN�fL��V�Gk�#��hw�T�ś�n�Ec���2��y7I�f)YY//�|�$+'�.)fs�EA�֖�X�\��������i^������36V�M���:��<����V���;/ K�+s&��]�8y�Y�z�^�����)�bƠ����M�6V�\_!r����b�r��I�z�a|ﻸx�T���J�u?q��uN[e9�����N��SWt��/J"%Y�	�9�[����M:��dN��a�⪌z�
���g+�e?�שO�5���z�����[k����O��[�e��%���	�d��̩�0�C��>~o���M̵k��]��T�� o��o����u�nC1�U���sI����'����m��o���Ի�YތԔ��rb�mp6G�Z�w>�s��+�,��3��Z�9��G��ԋ�xkF���q�w���K�׷���Q!���x�m�fb��!�tF�*��S�|�_L`>���*���)b�a�s�lN1�Y��!��sǎqbc���z�����������	+.D鄡��'5��5�a�$��T�!m��aS��e���:��6�h�SzUM�?bp�8�?� �[�\�p��>�y2Sc����Yx�>66�q�p��ۤYFk��G$^����Q^��S,n�`w���X��d����s�ӃC�Vą��!Y�=~�?��'��>EeV+�]�H�j1��7���ػg���l�8���#����2N�L�ͳ�Y��NZ��8��˯c�g��	���� �b�x�QR���Bm�aÈ3/"����q��U�{����ԑ&�x����tΨ�l�ܤ�I�;L��n]������g��1|$Y���q�Y]R{�`y��w^�FP׆��.��=�v�����P�C�-���ƿ�*���t
B�,��Ӕ(�l�-��nr2��-�b��w���U�}�S�`�$x`���>���
���2�\f���2�My�~�ן�<��Ƽ�M��!�7�It��3&��9���h{;�a�b<��C���r��z|���a�X�(V���[�I��Hr6�a_��S���k_f����+_c��ϐ}���z����'�K����]l��=�(D��'��'��'���,����������v���+��{��sz�\f��>ky��3L9b3���O�؊C��CZ�{�o;bmo��ވ�����ሕۇ��ǲ�y��l���!ɵk��)��ɿ���7ѳ����t�>���+�����X_gZ��`9�n�>��j5Pf_THZ�v����;V���>��d�8�)3�ǹ���<{�@X^�̗I6֐�6Tٔ��]v&��v�A0Xr�]w��m��C�ͧ�B::�,/�;�S��پq���.�{y��2��ܿ�����E���+�9�,c|{Q��V9�Ν&�m,��<�_��ߠ�Z�!~�������M����tz\�xm�>x��+W�~��{�{�8Wo��o��N�/�	��x�Cf��.��>���S_#��YZ]�/R�V3�~��tyI�����gٸx�[���Z^!�t�I 	;=�ܰ��ܺ�M�,V������\�y�Pֈ�;�\%Uה���<�8�1���G߾Ҡ1����s�g?ɷ?�i���o�Њ"��֖�娻.��g�����y�o�Ë��/���}�ܷ�cuL�5k�	�%�wI��~+�����RԍV����h/2��.�r��<�l���%��B={�a]�MK��}����m�\S�y�HE���]�G�ù����>M/:Gq�$�O<���
�AjX[nc�y�O��Hr���?�iҴ$�����?|����w3/rn������m~�;�$�����>��~�ӛ=���$,Em|Yb
�L42�xi�wލL��0�P�@���N�Cأ�k#���[���,}�Q^���������uͦ��/Q���B������|+A�1Ѽ&��@�DQ����#�+'��v�����L=�L1T�N��sϿ�MB�a�Ry���V�Tq����v'{f��3���鷸�w�!!HA'�aH��.^�[ܼ�C]Yt'�.2y�1޾~��r����J`1tW_�b�֘��^a��oܺ��{.�9�A��.QΣ� �4)�I��bL�m1hu�=<�����	�|�i4�~�0�jΟ?O�����h�������$��S�w2=<�(�k%���rj���y��<����Ҭ���s����#��	����]%�JR��(�4'�Rt:Ż	EK�\������Y����5�tN���pqHu�|o�]������ҏ���������,f7�^�zӰ?�2�eMҘ��g\��5[ӕ!��E	I�(�}��JPǶ8���0�k���5t�=}6�A1�rK�Ƒ�$m�.�[��ϲ�k���P5�v�C� }	ޱ?��Dǣ���o?�V���T����wn󊮉���8?�������>�I6Xe�5fs���h#h�	�,Ŕ5IE/�:y�pi�0��N�V8!A�D�;C-�I+v�!�+y��/�x�eZ�S{CW���D�����۠#��q���!��E �qf���*�Ѝ�04å��I�#I|���`㞻��	Ei���0�~�g����_|�JJ'#
c)��N�����|��x�����c��r��;�y�F�}�(��{�Foj�^����t�֖��&��@7��ΰ�1s���U�������~>���+'�y���ٸ�4�*��w��O��oq��y^x�e�()�'	ݵ�^�±�w����<}�7^���ub}�|I���J����O��o��%�q������o^��{���믓"��LNYW���|��1>�(����V����g3�o�e��mm	��5�a**��AH7�0�o3�q������ݥe^���y��� Q���)������:���(�q� �;��+_�:u�Jn^��"[���S���� CAi�I��R(Wsbا6�*�U�4�G�X�w�y�9قB(F阪���`���|�*�kj�M�I�����^�����S�]�	�=��6�*J�J���gv�`���a�j�.b�1�NB6Q
O�.y�9�����+<�Q�\Y��6��Z1��H%ą�S���Q��u���p�����"��p!�R��p��;RI�i�$$�T�`]t��gW��������0�)�&����B(��P��(UBZYҬdieH4 8����\�q���m�߷�����X��BV���>�g�gooĻ?x���:�m���{����g����=-��4�X,fl�}���e�:��o<���;���l'�$�xL-�_���/��9�Ɲw���*g��������W��<�єi�#�bv�/�tA�6���w���ZZgϤL˂�8EȊ�	a���&���
����أ<q�#�w�<��~�2��!�ǂgk�ׯ���Ǟ@-�Nr��%dV�j��B�NX>�A^&�a�ng	�84�&P�����ы�n
u�`2���~?L�c��J�H�`.Y��� ��␓�9"	�%'���2U0�Z�F���T���"G�!����Ֆ̲�d�E4���]A7Ӫ֢S,8��^��d�`6c6| ��/=K��$.��l�9tܿv�W��3���7�Y�68Q!���'E]���z�� �@�U+e�k��1z>�����b�fT���hE�2�,uZt;��-��	E�49���=�&C,mt�L�^%�(�#h���e"٧��6��� �����N8hintIҢ�����=#8�Κ�~��r��Q�٣��v���PA�R���3̶��E�1f+��U;�޽;+tK�VD��6����I6A���16>�؈d�|�H�c�:��Խ{�Ωr��k�<��C�����U�z�UUk��7����i��n����C: �$��<~���c�_�܃5jg��3u8��	w^x�5���R�MJcg��+/���������(�^y���3��2r��e&�:��A�����7���@M&����8�;5G{�M��M�Bp�p�mo1�sJ� ���/�@˚2�{�Yr�K���*�����4�IxE��fN:�7.2{�I����5��_�ƍ���{�z�,��1��a�D�3��`�0��̧i_y��θ�}�'^�2�w�����+�6e���f��ka=��ŗ��4�מ��ͧ��W�[W���d'Kػ5�m��AHz���dw݅s�fS���z�F�e
Җd\{���h����_��.y�b��W2��qiCse#��[C^y-�'/��>Ĕ'�ěq�Gp����'�J�E�x8�6�@�F��̔�6=ܠ�T��5�����p7w�_��ʸ��"mҜ;B>ڇ��Lp�2^k7�aa3�f�~��G�#'2�70� qz��?���F�E�y�R�u	R�H���j��&�~���2����k�H]��!�F�u V�����1F�d�2�>�Sa��AjJ�@�H2%B��ДiF�eTyN�s���\n��i�9�C6��B��¥@�������
G�V	��8�I���tJ�բ�I~���/4�+��~8����TdIB�g8��g$�o2}�U�����oq��_���+�.\���i�d ��*����[����מ�}�E�>�W\���(.�L;�����`ڔ�Z�B�Ez��_|��+̾�$���o���"�t�Qf�{�����ҴW��ސ�/=�z��W_�{���R]�M��XB0�JАf�6sӒ�k��������>��g���O}����4g)mǣJr4&E�0>�N�q�޳�3{�y�3��������	����*����� ��r�I���c����y�����l�+E�wq��db~�4(�M��EwT'd�aH�d�Ki�a98�K*``����~cFY�f��$	V�@�b(���R 1@ο�J�6j8dɘ��K3��U%u��w4��6��Ϣ6hU9i�'+v �	`�h� O
��Ȓ��6 YJAfq���*E2�#�y����,�Z:�ל�������¯\�Dg�p��DH��`6Si��&Y^`���a�0@��R�deNfdTfIf��t�r5UhS�	�LA(JQ�)0T����*qp��G���w��<��D��w�RNv	]����.��:��P]����:U���lJ�f�y��v�f?f��g���?����"��+,>K�����^kb��B���>��>��K��o�0��9�����Q��)��疏�2��?M��/}�3ȗ/�M�[�����@HL� `I}}�������`���м�O��¯��$�+
�p�!���ߋ0^�F��˸O]anc�Ry�/-˒N#��XH`�9:��5��/P=�
��-ڣ�9l��$p*QY"�ROp�������㽺Ak?����n�`��1&e�b�[{�7w0_���pg�G{VbF�t���!����uQA���wi�.�-u��m�Jgu{�����?�L��aZ��Ժm�F� L�3�8��]`�b�b�ϰ��EXi�S����r4@OGX��QD�M��m@Z%h�A{:��d%-ˤ�����i��&l8;Ø$�Q\�<H\��+͐���'����-���oDK�j4m*�d\���m���"�SF��BV#�t�*������1O0n��Z�aڔь�קY�&�Y���b�6~�Į�0�T-
�$�9G)LU����5�*���k�����'��%�����u�T��=���=E�J���\��Lf��o���t��!q�:vqȶy��yO��Rr$*x}w��ЧL6J�CR�T1�-���<�9�9j٬:vR��®�\��Q�ɤ�:��PUN+t	(0&3la�t�4�H���>�a��۱A*,[�P)yK�`�@�đ��C(�2fT�T�En��ml���,��BN"����֩��vhk�X���(|I��8�1�x1�'�٠�M�]Ӷh���۴�5:Kk�C���n���3��P�qj!�N��7c#�XhP�S|s!N�B�,E�`�,v�N���an�Ԁe l[�CZk3���I�g�)��:L�L}�i�r��89+YL5��Q�k�P�]AU�h���h�h_!�T.T�f?���3a���aq��q��G%*"H�t�F�c��K8�u1}�m�+�-0�PL�y�� ��
-X������K��v��7Ü��2#����[����s�q:"H
�8"1v�3t0M���A��˒�ᙊV]RM��1$�&���)��C�E�v٧���N������O!�a"����08��,QB3��`��^=�\��H���'��!�k�qR�t�$�
��%h{���(��^�ƌ�Ic��H��	^#�
}*���ܔB�pM6�{��8����ɪ��Z���\�8�u
�P�G��0VW-#�u��˄�������iZ�u���s��hx�(� X�`v;�N�x��c[��A��dya���"�����<��.sw�8��\m[�~h+t@h��{�ss]YP��pϬP;���֦yr�ŻO�=sx����9w�,��9<i ���'�[�Y��~f������Zj�xh�?� kGa���ìӶ�\����"�`:LL�hR��A��BLe�J�mb:uªN=lP���F�j�0��)&E%P�����ĔR;P9Pؠte��a�&�8��k�HsEX[��k��K'�����q�2<��8A*�1;��}7��{�$ȝ�
a����G�����p5X���;'H-EE6��]9ʆ�Xy˻0WO3�w�/n��6E���p�p��[A��5�
�x~s��]��Gb����r��#�z�R����tERdh!������lF�2J�(EEj)��`���j��P���V����3��0�o��@�����!:nJ��h�T�p͂���[�l��L��6��.gO���]��b4|f�D8&fˣ���@�J��kղ�}�6	:5����vCZ��F�c�>�*����:~萫�</)=��,"�5u�gSqQ�1��/��9Ґ8�G!���̤��Mlϧ�� -����|j���_�Q&���F+�Ia�C��C�=r�D�J+ꁋ�A2��l�qHm�\�v���2�`9�u���$����Ėi�H����,�����{���e� Z�:�n[HL!�9߬�=�Ӵ��B��jz�`'���ǘ���e���4e���T�f�1*�T��t�)5�f]kv<�ݺǶo���LIZk�]�F�8h|yM��g(m��;r��5,�Qa���ؔ>7�r�Q�0�*���<7���lTw����y��e��ڰ`c�����
(M�m��\ff����m�k1J
��2��s$+Tgf�,��cty��wq��]�<r�����<~/�]�X���º���j+lV#�ɝ�2dTٌ�K�������U�Q���o�zuҰEϴX/Kz�M*<�<@Xmt�� 'SX �c����� L�3;3�Gi��:|��z�<-Ѳ �2,�&�2<��w�ԃ^�-�ب(����J�6+�T�vq�tc��
%+���6��C%�퐪�J	L��ւ&����OjDZ�f��N�,�KJ��:%*�g}�-pM��d��Si#�&��Ɗ$�qHa{�����4�Xi�cT&����OP����iJ�Ԑ���~��Gʹ	
9J11)�G4�"f�+�����:�6�c�-A^Z���i^�*M՛bg �
׵�~&�q�M�Ճ�1�~���(e0��<u�|�C�7��6��2M�	A�<�MǸzF��@���^B1T��w>���^��������%xכ���QZo}���?��M��~{��a���<���a��v��f����5�#1:��9n�������<�Y�r��t������z�������w|?���c��s�O�,o�����!�{��<�w~�=-������������\�aj�2w�7���cw7����.]�l���>���eN?�������f��v��q=\aôiL"Z˫��>2�)u���c9����|h�*�р�Z��~��P�X��]�ѶEc�F�ݧ�5(̂O����=ˢo��%vR�/�A�?�^&���?��4��*���Z�S���)��Ya�e�8��L�&� � O&�W�^9�%8B�\�[8EA�V�� ��X�D��QP�
a�� �*�
� )Ll���9^Ybz>�ل��23 �*j�O���l����I�|���U��9q�~���c�?�eYԄ�5���ܒ䕦^��5�4|bYb�2��=������O��a��A�n�IgY ������@�fh!�F{۔��Qh]1��y`#*�IN��<%��TŊ� k;LU�.3X:��2���:v�a�%������`u�͛��:�{�������Y�"f�a�P��.m������<N�wp�?�G��&��ʔH�c��W��_�U��`0ؤ�6�l��.�<���ցU�(*�q�ؔ���#�B�Bq�Q#15j�ե�=���یT��bj/�6'4�	*�#��۹�ů���*}��L%$�7Ur6�=2V��:����ͥ�|�s����xB{:厈�>�3ب�ukBgi��x�ki
��r�L�ȰE�T8���$NS�,'��0�f:E�
ג�q������c��Tq ��=��vjPK4���ws��IFϽ�_�;�ȩ����h��'y�?�4����1� ����8�m�S� �,J�g`����;�;��~_A�Ğ��aQ��� L�a�X�s0��A[
�5�-�^Bc:V�i��^���[��8��wq���D5�k_}���]z���u��7���k���6]B�N�̝����W�엞�z����w�&3���gM��gϱ)L��gR&D��pu���}�b�"���_�C��ַ��q��q���
q���u��0ÂF���5�:uUT\���D�7	Z5<KPV9�
�2H������D86E��T�y�M���0�R��0�28��A�ຒ��N�B���sO1���S��%�?�Z.�e�%1��4g����
a�$n�^����.V������`�tss����iɥ�M�O� �KB�&�Rr���C��\Q�
�0(ER��4
�n�dbh�Mћb[y���,b��?��?@3�Q�{�[&����W^�'~��Н.bkU� ��8��Ђ���9����җ>ˍ���|��ϛ���i�,�=���4��3O>O�k +���u�b��I�hX.f�)��p�Ѵbcg���hϠ��������/_��K����>���wqrn��W������6���Hr�B#��@e`�5��<s���_�1��}���_b��O}�����h�3	�,B���k �-4RV��$M0�_�E�[�,p�`z �I�4���tqp��B��2�(�Xh\�³]� ��ٯR/`��q>���� ǽ�x��X������mN��z����
���Gx�(�4����~'7�w����;���d���[�i�c�(]�u������?�ܹ9FZq��7���-�������(V���.,�w��M:k�(�e�������3\������q��g"�F���d��h���,׷p=�Z���MǠ�i��ql�
� ��1��1�u�\��Q�-԰�9à��O����c��gmw��q�� ��+d%�*�J[��B�vY����~�r�sO��Sw�O���C�����?�����Sw�z�����Wģ�2ͨ�.R|,t^�J� ��^�^�QBZ��r�D1�����paZ\���lX����]�Y8v�3�����Y�n8`y^@���f7 ��Ԅ\su�Gv�	��K�?y��9^��W���>�~���}�}�J�E���i�|}�t�0�� �)�=#Iv����S9����r�g>	�LL��K��!�Ma�,�9����m��7?Hr������ǣ��6�w�l���E�"Q�J
����BnX�}ɊۤHBiӵlj��ƭ-��1��03�k��P(�c�g�l��`o4eTU$֌ܘQZ9�[;��R�LMbjҬ��518��e����EIPT�y��2��iBo���`�t6㓿�{=��C��dܿ�p���~臿�8���&�d�p{���>[�!z�Ea9�K��%Mx��GI���=��We���-�ܸ���,z-����C&��഻�v���?��A@Z	ƓI�0�bVN#�*���S?�����E�no�M�����Wkj��S�Qhɤ�qs���`���O��3��'�M�o�`�aG�#V��F3˱�
k��
+��a��@M�D��˰L�,E�Q���6�,�5+�2��9B'� �t8$,�Zt�,7Ln�)?�s?�����_��S��MI�(��f-@�M=��F�9�-�4j�RL�I��j̰��'ϑ�	����3Fٌ����'��?��?dcw���2Fu*��yI�����M3�7IB)LAj	����<�frZ��&�$e0Q0�N��'��i�RoyIE�Q2�1��&.2q)J�Rb��D�F�vh�.�%�Y�ȍ'4)���hȝ�M�y��<���|���+~�?�_���eR;g�-�$iES(�|Jˆfh`5��fkJ�NY|U-H�A�.�?����<��}����h�	���� I�����w/3�{�O9-��ꍱ�nb��q��8\1�	2�GߺLr�E��/^z����?Gv��D�/Sv(��(��Z��.f7�?���������?ae�ςo��Ǒ/]$��x�![�n���i����`����!;����w��c�������c��������`/�D�y���Y��.3ڿ���'���_��O���EQ���� �Q��	ލ�L�/�>�jA�J`�퍩G>.������_d�dE;���49Q¡xƉ,洨���Ɛ3,S�$FS`6�(�f<@�ߦ�8�[��m��8�g��x��!����ʧ�W��[�x�b��B�3����y��P��Ɯ�����j�����|�'~�ct�.o������JTB"E�a�h�����7��e%n̀(Q�'0�}�iY�7����ת��#���Ͽ�;���$���h]�LM�H�(s�M	2�1�ϘN�f84R	E)���`����E	�n�A��ٌ��dae���]��{?�~f��m����e(� �b�bJa����TB��H�>�g�f��,M@�r�<�͏��Ck�i�:��'1s�4ϩ��9k��\V��,�k:�X��)McF��i��2e��S�s�{�(k�:Qr��N7���_dAT�-�N��*�isb~�{O�E�pp���Ԙ�e�G���9��-x>�N��n���偻�r��<t��{������>���Zۣ@�H����n޹Ē���g���q����,������Gk�R�&�?��\��Y�<r��p������.�;�RP�3-���lM��Q��O>������<���82�1�Ƴm�y��#,�B�C�DX�ﹴ\��Km�Y��qצMX�$��m�;x�>DxY=L�r�x�A���h�,Ԛ��j_Z��m�߲�l�w��ݚ�Z�e��2_3hV1�rF-�Q�f��9�%�}���u�� �ױۨ�;��}���;���_�VԦ}��w0k5��;���>�"���U��m8��[�YFEA��F#�Q����d�/-�J0�*αJ�p�ŕF���/-!*�rؤ���P
U���6��&�
�<�<�|�JCUQ�
Y
�J��+*�7��?ў?��}&Q�ի��B�����o`Y&���1���('�)�1"SJ7#A�
�P�f����C��t�l�F��}�>ȑC�0��Rx.\�L;lb&�ېXYFk��'C��	��=E����n6Ƙn�dcԣ�M��S��?K1'c�q;��L&���Rf��2E�V�H! ��qL�<#��B	XXYů����!A%�E�RB($�2M��?�x���y-�ۯ>Ou�_A��)�?�U��>K���*	k2��k6��*{����s���a7��>Cv��ŀ�����C;7G	7�}����ncC.>�)��g����>�ISs��_���F�1����	j6��ʌ�_"0s��d�_%�Sj��R"ΰ��Ʉ��Id�a���a
Qh�$CT�����q�d�0�N�Ɩ
���;�PUb
[�	H�*#���"�*Ǟ�b�3�x�̦X*�1�1F^@R��*\�K LHd�Ցd�.���1UQ6;0{
a�5�7�4��T� ���Jꅦ#L�l�m����Q�eJ�Ͻ�/?�<�(�(*����ݍm�f���a��
�5�a�@M)��&��Ł�ğ��u��=�lL�6F7o 㘤��S��4����`���N9�U�a�sx�<V�
�"��L�q�2mQ�-�
�����GZ�ڡ�{{#��3ܠ�eϓ�&{;^x�kx�O}��r� 3S�FD�Ed�aF��@*W�x��5����O������<��DO��Gj2BD�d��h���@2%��cPIA�+,]�&����8����aw�ǳ�Zae*K	�3)��G�HU�n�(��wi_�M���?��`D7*77e���5r��Ըp�6[�n�Li�-5eqo�ۏ�5��שm^����Ԅ,��%ҳɷ�鎦x/}��i�o�j�����2z�	j;;��>z<C�%ZV�z������X�,x�N<ĸ����*bD�`�RK�8�_~����
OWEIXT�Z 7���)����=�y��&e��r�1�$�sv����W.VF	���Ķ �b��9�)�d�t�U�.���)�v�t�MYe�瑷��4O�E3���>Kok�L��l1�����0p]Ƕ�M/�Jc)p�
;/�Ī@&A��"�=�o��ۿ�����}�O����	Y:c�����iE����P)4ij0DE)���>� �����xx�C���F�?��?���<�����
�B�aǷ���I2��sJ+afD����)I�)J�ECp�]H�_��'y��'��ܦ�I��4+�-��w�����BQB��
O���Al�v�6F�e�'��&p�%�MNNP7p��X�EO�\��fMH���.PRb4M���u$ZW�:�PŁXHk�7��z��0MME����@A�P�]�B���[����>:��-�ӶV�:ua��`g)�"��g��UZu��lv ?�g�YL#�P+b�d�J��$�I���*g�~�Wo\�c_�6�^�Q�,f���N&TI²)hN',+��&w�x�/s��u�\|�"�R�S�*'�Nq�I �*(�1V%�Gcn������p�5f�,�M:�Em0N7��M�b�2ۅt���6�3���Y�C�	�Qe;�.�h�OQeJ%@�A4���uP�(���tJU�(�	�*�l�1�)�2�����+���+ĳ�̴������{S����lli�+ Or���"+H�5H�{�M�-C���m��q3 �MT�%�iQ�ygD?�a�9���+��\� ����$L�1fQ� qP��@���,Cq�y�M5�a<����_ᩧ�e؟������an�٥U_F�&�j`��@ ]��2G����+*,Cc���bY�i���	�@+A����K/��?dkg�J�����C�GV����f3ʼ@j�,�1d� �Cya�d�i�p�2e�b��&�I�x�����a�1P�If�Ob��ǹc�Q��W�K��lL:3��g3fi�p3N�L���7��#K�Y�0���S&є�hB?���L�cF�1�x��n�o���2ݺ͸���q���.{��l��0����b��G��O��ϣ��c>�hLThi�2�����	��(C�����$�}�����݌�C��w���Ӕ��m��)��-d1��`8���ǑC+�;��:&��Mv��������&�=vz{v{��O&؎�m�����`�A�pV0�sF��^oLowʬ1%�&	�Q�r�M�fT�L�����2A\�̴$*M2m1�J��!+\��#�L�M�8��hd2�BⲂ�%�;�_߂I
QFV*��.�ɄKW��4w��CǑ�&+�"m�4�iS�
C��B�����e���q\�i���J�g��������m��o�\�g2A��9M� �ImE��ɋ�AF��%��S���AB)5ɭK�:{�;��ܹ|��W��as�=����4��FK6Y�T���� ������Z��@jUTh]b逼�q�6y�#�.~}��#�X=� ������8{��x�_�/��WX�����ܼ�Ε�{\��˕[;\X����=�^p�ʈ+��ܸ6�ƭW��ruȵ�#nݞq�攋�G�z}̝͔��>Ǘ��=�bH�v%�����׶�}�
�n��ՋW�tc��7�\�����VU�G_�+�8�Z�׮���[\������n�s��-n_[g��%d�������w���[$��Ϲ��5p{o�˽Mv�)�;SF7w(z�ϙc��7[��۽Wo��ܙq{sƝA���+76����h���E��
!4�|��|cg�������}v�F��ﲳ3dc��p6ciy��_Ze�f���Q��0c}�s}�5��&�)�<�ql�:|���;G$s�F�31Xl�6{9�0�ZL�Y�:��2i����pk��Ul�3��Elr�{�;�%�;%{}����(6�
z=�``��{���7Sn^O��
*x��M����6o}�],-�3�i/�x�{����2�0)�0)�"�s�Q�x2��3��Y�Q9���V��8��͘��&����o��d�۰9v�,>���;h4�iBa�.��8�I)<��"¶��P����K��_���@�R�]"&�tj/��{u��d�5�@��9�`3�]����\�{�W�>��[����Ý�w�S�ј�~�t<"��{��a�d<��g�z����2���h..p��謮�|�8�=��	� �U[eRT������5H��m�`��.���0��N/S,���>iå��;>�\�P�Z�.��G�Z��AͰ9�����c,�����R*��	�BZ>�|@Ԁ)��d�+/}�8)�m�m�FH�؂ɜC�uI]�����C.�z�?���6<r����0�T�&q=d�A�Tcڬ�C��D�!ZZ�l��l�#���C���3�C��ZE�$�p���sױ�t���u�c�y�À�7��z0�KJǦ՝���s��)�mF>$-�"��W氏,c�CT��Ա��f�����-<�Ƈ���
��IҲ)� 
Q��:U( �?��]gV��AV��N6��Cֶ(���9�y�ِ��$,����ω���+�9%S;cd�L݂$(1�c��D�nn./p��-.��_�{�y�u����s�ɤ��p����\�y�k7.�q���6o^��q���:��7�n9	�7�^��H'ěw`s��Ɛ�[=��Ɯ��;̔�g��������M����O����o �89��P����7]:ƿ���a���)���y�t�����5kl|�E&q��O?I��x׶i��c�f3�9�i�y�.�UP�3:���8�1bNz8��x����?LF��.��>�p�=R�&��a4�����h'SFW_cr���_��3_��4O=���Y��*ݰ�Ө���jsԂ&CCS8>u���ݚ�l���M�v��F�!f��vl�f��qAq��R���[�z#���<��2q�h���V1u�F�ۧ�_�[=���.�n3�L������k7�?i�8^�DJ����6}�����8��r��5�&�i`X.��F�I��yeg�i�A��;�(Ҝ��6y�cy!�S�ku�]֨9s�lI�p���ȕh���&�t��Fߩ�������h��:E����km��UnolP���W��MYHæ1�@�;ʢGA�0ǬQ�^;���].]��hoH��A��з��K,%c�#_X n70���m�s�Ý�v���I���
�h���Lh*O�=��<�Ț�F{�"?������ܼ~��������k�W\��
��u��[�7nSh��?B�VUѐ�Lq˜
�Hi�
;IpuJ;/h%^���lV�ؖ�3*,�ba�Ik���]�|峟����l=w�������Gx���Ï}+��=�\j�ۜ��;����c����M�������?gv�w���c������O�Ο�!���_�U��{Xkm���ocgw�O}����.�y���3�S��#��ID��ma �KM5JжEbd�Kki���aJja�t�]�ǒ�<�@W���F��&wx��)N�C���_��e��V.��PH�N�����Ӟk�F9�k�E�q]�J��Y�Z��k7ɖ��xCc��{���̼���[��v�,�?��\^`r}����|���<�v�"������Ԧc�I�ͺ�]�$gk�Ky���6��!L���)�_�S����J�L,�[Rq�,H�:T�p�KL�#��6��Gt�<� �9��\���;�ˇ���UF��݋_���;�ш�'��G�&SY���J��{_��d�����UN�Nm��M�b�+V+�W�Ʊ�\��z�Vg����_����_�kYF��+�
����a��t�9I^8X����1��w�a`mm���2D1E���=,�!ȳ����8���-�R!M	��R9���������쫏�l���,b��e�Whnm�2�R���1̪�څW���������)D��S�8��k�r�8'���ɐ�'��B�~�8{��3���_���%��Ab�� �����$����a��c�2Wz��~��Q� �NM%�Wy������o�a�~�?���>HdH�Μ����?����}�=İ?�t$�ş�_��?"� ���u���u�f��.�x�h�~L�f8�Oj�{�y�$�R�&A�I��&j����[��,����/�Y-^��_e��WY������I,�;��\a������z�C^h�TT��1s�����vWX~��qa����Nݜgs��c����W.`�\c��WI��ޙ���DS�b�uQE���.K���ְ���,�O-5��L&}8��F��Yc�[���Cd�����i�&xqL���W�}?�A���gx��>�Kǐ��7���cg0w{��oR�}�&��a?�x���cO�H��a^h��M�?���S_Ùi�c�r��ш��9�挛Q��S'ʇ����6���[��寳6�vhϯ"�\?��p��:j�R)��p�X��=�`U	�ן�v�25ϤWV��{��z�sqg�v'����,�?�=��g~��n2��[H"�n�P�>E��	�E�]	jN@��,�iӓ�q�&gq��V��Kd��+F�&K*T���v���Gd�&�c,!0˒r�g�ߥ&���$FN�XZ��v�;̨�Ӕ���1+XZ\ĩ׸���(����È��Q:����Q�.��~�U��vج����x���$� ��HOL07�������eꝄF�i�2�}/��߸�
�֎Q���ҚH��k����yu��;�ϟ��M���ʝ-�Ò*�
mC�	�Q�a� Jʲ@K��a��J"����VG��y�*%u�`xQȨ�'�,�\�i�������\+T�&�"j�FG)�c���������ɿ�*O<�y���^�������w�����w������gs�e��������o���!/~�<m2 F�&oz�����!>���GM��:����o��sڧ��_�/o�RU�ؗ����x��o����B'S�Z��d������������'���T�������?��h%��_�+��vhT��]��>��؜F�����j�y�����?����#�ʏ�0�tJ3�P�[��x������G���Dۅ������=�������Ѫ�l���*o���_|�K��寳�7�̃g���>�wy�����G~��"a��E�P=�c��'�3�����&B��#Iwm�7�����㳿�+X_�y�n�&�v@j�X!�0NJ|l�"�
0�6`��m��X�^���	F��d0%6!��� πz��VD{~�����P(E����B`HC�HK��h	����WV��o��	�� S��$��I3�X�ܹ{H�lp��8(����#�Ĕb��H�n�Z��8s�G�C�������yN�eԶ�i\���fD��U��^�4����s(���ܡy�ޥWytq�CB�Ѧ���?�S��f�E�*�eNf�T��4-�Y
�ԋ�Z��d��H���U�gշY2:yN�,8�4��VǴM[(�$&�\�ZI�*�,�*Jj�@`"�!��Y������=�}/�����V�׽�Mt�VxǷ���IX�(��vX��4W����i�,q���9�^Z�E�t)���LTL�Qgg�M������X=���'iYa���9s�������w�;�P:'���񄉚.v@Y;�Q)|Ϧ�ip��]�ͦ$�� ��Q!WЬ�;�>s��Y=����5���X�;��r��t�{�ַ�9u�çOq��=,����"A�ͻ��1:.S��}Lz����S�}��=}��ㇹ���!�y��x���K�
p�I��[XA��Y9{w���Sg9�t�������.���w�k�=�E�>R@�s�*G{���5)bPI��X��8ؖ�V�*���܅6YoJӂ7`ٗ,�rR���&g���K�x"�&
ֺM!�c���{0Y�X���>�Ɉ*�p,�mj��6��5D6���9��j6�.��1�c>�y	+cX��`��lȲN��$�H`J+����O~ت*�阍g��u� rp'��э9�MW_f�ob ^�0�8�t�C�Eʼ"*J:���5�z�a�1�%��33�e�UE�ڣY��:�4��
�u�EY؆�LK,	�oaX&R	��²4�a�&�	n �ɾ����m[�<���&�.&���)�N
Z�?@x�4���`��*^r��Y�z�,�Nx��� �+UT��X[��[e��)N9A>My�w~'GO������+�|/I�z{��m"!��[���as0$)
�0��|�wq��S��7^x�ѵ��M��{�v��Q��s?�����"g��Žox�C�N37_ÊǼ��O��Kr2�jJ��Y{���L���%����c��X��\��ؼ���P�D��;��"X��>q���az�1�N��̩s|�?H�S,��y����(&��s��)�����v��}�Z��~�����g��f��Y���?N�$XYEV)�z��c����ۛ��>����b��������OF�h�x퐪�	�9\��d�u��!-aix��Ƕ�8�e6��F��!q�P�&[��ceH�����bJh�bVD̊�VG8i�8�BP�����kӵ\Z+]�"%R1�'�!�<a��Bͯ0Jvp[]q�����d�5������;�y����0~�C?�a���w��˻�d��$��%�;Ɩ���Oi����xJ������p���:z�#_�Rf	v�NNFlHD`���
�QfX�$p,Ӄ��*�� K���R0+01���Ԓx��5�Rb�]��EA�y�|�W�Hl�РR�cɊ��(<��
�����yR��zca��o};[y��o_���㜺�.�������l>�"7q�y�(|���ì�u�g_|��������j5y���QN������e�(�hV �Ia0w�8ۣ�C'O��7����{��7�y��k8�OK�k]R�2�|j�O��/s���t�$ͣ������?�K�K��F�v1���r��Ԃ&'�=���G�o��v��9���İ �f)�����WorsoB���o|u� �]���O�����ͨ&�,#�*��}v���ė�|��8vt�_�2����������6���w�-�_������O��6��ef׮r��_������5���RIj�CaI&�i(�J1]���(tA.�J����1e�jm����
H����`Gkl�G�M���>�_�v0d�i�N�l@ea
�x���!S!PINm&pL��o|�mSP����\T� �kL�:Dz�F��쭓����������dp������x�ko}µѤ�R���5���_�ޗ���dJ��R1�0�����Zs(��B:�]{�sG�A�bl%��H����FJr9�@��r<Bᣊi��y�\0�E$e��8 ]gY�4��P()(���i����Qm��[��v(ҜX1���\,[�%	��+E�4�
,Cj��$J�X�b4L(O�B�� ��g��Wo^��Ջ��p�_�<�>�	��{X��:�H�ǖx��=��#l��bo����"O��/��U$�q��z�"��X{�[Yy�Y������u�z�����=��7������ot�Or��g�o6x�~��ӇQ���,�$��g?����XOp��qL��PT5����~�;y�m�rsڧ�i��F����?�=把��jQ�p��8|������C�g��h;L�x�K_���¼s��m��m�A��R���H�9���<�j��O����
/}��0���;���3����G��&��>��NZ6��:�x�����$�p�����M̹�4ϱд2�ĉH�� �a�����)��$����g]���1�Cm"�`��Ԭ���F���[wH5$i��M�Y.M�
��0�I�&��M�xJQ�hUJ���{�}�'Y؜2��F�7��wr�٫�q�������)3�����w�{���W1Ҕ����It���MJ1b�5���_f����6y��>��[Cy#�����%-,�}�~nಾ~����r��	��&�e��+ϣ0hu���O�Kb��M�4�^%4�*�'I��y�EJ�w9s�8�����n50\,��	b�z�������s�^δ��U�z%Ȅa�Z�BH�*GW��U�+��`i�9��h~����4�D  ��IDATLcqò�m���mn<�$�,������׹{�Tct��m[������`�*v}�9���W���M	f9^Ӈ�c��V��S�{�y��E�f���ړOc��(���_��Z��J��6;� _Z`�����7vb&/�k�?�,�<G_����a� #@ܿ4�О	��3v-�'s��o&/s��^��3/�O�xq�lk�r�I�Ø?�{�8��c��V��5^~�Y����iA������t�&�)N��N�Ѿ�n�F�晓X���r��5���Ʉݫ�ӵa�u��d��}�iw	��i����4�w�&;W_��ol���ߡ)l&y��IB�Fٛ���{�g�� �)s�� �^�>�](f�]_`�=�ͣ��_�+a�وX��Nڋx���_�-�ˋ�$��$)F	�eaYeYRVm��i�g�ED]	��]:�:��Q&%YC�S�9�8���vC�M��{���n����������?�he�ʑC���~
ݭ#f�JKb��k<�s?����=������U�oE=��]�w}�n�����絗_c��I�<M�-����zj��&Y���@b�S�_�$���*�J�1�rni���ԥ�/<��²=6�nr��x�:�������O��G�S���sI���%n�F��24��ҤP�A�V)0Ra*��6Ci0�[���(iPi��AMU�qL��qC��C���eJ$2]%-R,�@�� t)�����"��Cc�ݐ8��k�lo��w)�!e����t�e��)U!�uZ��$"���	q�%Zn�d1^�@h�]�QB��I�j�0@��A�����8KT���!���KJb�gLv7�dI0�A�$E�ޠ�ў�[Y���FH^$8�kkD�vL�Ё�p}�tF2��ՠ�r�ҵ�}�JWhUQm��ْIt�8m� sH�`/�质<l�
�t��Ċ�:X�#�ߴ��
<��J\�B���@3b9PT�I��Z�������>�����/3�����d�1*�9�K昭�A��eE4���ϨM-l *(�� �YtSaK�M���SUF��l��͙v���'?����o
�¦��oma�/���������E������A�����_�t�C�f�V�8�����05k�G��?����.�O~��_�׬��u(@"Q��o��W��_�ʓة���2����QZ.5�EX�YU���5$n^��F9��TiU`xI�	D�B����#D�>��E�VQ���8Ng��o��o�y����x���2'�53�2�QPY�݁\�誢
*��H�0E�V�e
?0Kc��1��eyx��LW�"G�	�=dpJ��#ju�bw����x�,2�]2.��Vx�GUoa��T��(�qI��T�X�TUE�f��`�5O}a��$AePsl��yNYf�d��5�
H*)EEe(̖K��DUNUiD!i����Ӷ�6-�$�
�0��lK0��}˒̲	��a�X��j�*�(CM��`g䶂��V�J*��	��X&�%i�`�wю����(�y��H!0��(���#|R78Pl�3[�tC���$I	r�%��R!�Ĩ�5��Z!�FX��S*��"^q:|��_��Gy��>ŷ�����ރrltQa�f|�W��o���ޔ
�3�Z�� �E\ddQ��{���id�E������*Ƣ@�\������ݼ�]'N�}��wY=���b���pȕ��c��͟�����}�'~�07p��Y���
l�����0T��.�?�7�|�wђ_��?���<�&�#G�q���7v�u���=n�v�Z!��O���:&�M�d"#.��ў�4�՘%]CT��!d9�mC���x������E	�<�&�>xۗ^��K_����#��*ӗ�a��qbM�0Y6+���Tt��mL�74MU�5$M*�@Met����Y.5�Z�&���̥	�`���!kńecJ�G�Y9K����L�,%U�i4V��G���36J2)iaa� 7t�-�*�R4���X�d��9,z>�`Jj����,D^ �� �Shϡ�I˜Ri\e�(���0M���ԃ��R�굀Z��������թlI��it�Ԃ&��R�}�5�n�A��B����:$&�l��qq=��\�V���ai���ph/ͣ��E�@8>үQց���<�M�VР�x4l�s������a�UPB��y�#,�4H�UV8���dE�h8%���Ӝy�1��������=Ǝ	~}������'���^f� )�
�%�e���DEeJ��C���ǑX��eJ�W��[Ǧ=�a1�q��k�Z2�p�=�x�co�-oz�N+Ĩ50�i���e���"���a���Y���/49����])�H��(���@XP)Ʒ^�3g����D��xʯ��_�/��?��>΍���a�6����J]�LV��4ҵ��SbyU����J�|4BGS���gX�v�z<��S|�ӟAK�nը�q��'OQj�	�l��$bioFs< ��iL�4f=Z�1�� ��E0ޥ6ڣ5�M�,$��L�T����w�7����޹L}�2��k��l�F}�5�[���a�]&ۻ�	����Df>��c��[��Jq���/K��U7鸊5���|�NQ��%�M��5�E�Dc��-���%K�(a�qX5�oq4�8�q���r<t8+4��p��8m���<�C�Ê�Y��f٬8��1�`�T�����X05�*�Iμg��9,�k�����9N��.8��Os֪�%Y��][�J�tJ����'�D�SV�)kքSA�!=�p�r�4Y�֒�ê`-pYuL�Z6���ZrXV����/��p&08b��
��-η<�d�\:刬����Y�e�ɂ�p����S�'{��!_��'i��=p�K��Q�`kJ��~�,�(sh��̵�TEA�&������͍�\ؾ��d�礻�:|���pC��Jy��'8y��{�a�Ҡ%��:�>%+����H!�t�KY`]��g~�ǹ��<'���{N:9·�;�?�V�~�׾�<�N���_�
^�ƒ�@Z(��%\�Jc��`��Z"��4�q�65���M6�#���dJ+4x������ɔL�$�͇���~�S�.|����V?�g\����mN��.�Rx�da꠽J'�
�q��	@�9e�1��E[�:ÔvU26gd��k:1�p�W>X�Ԉ����I�f����&8EY:�a��i�$&At��������
G��IC]Y�YDIR!ȳ)�Q�9V8�`֜�`BU&dQ�v�TT����3��f1�N(m���kژ�&KS*�!<��
��!��e�U��X:�H@��*�,]��H<��bfml��>I�Ӄ�}i�%`ր��������*��r���C�PP96�̱�ب�� �5����ir0&�*���~�;x�#��W����Y�ܿ����#��~�?��W_�G��w��J�����PR ��lL�ԚM�v�*���_X`��C
J�t��,6Z���d>���r�����R��q��v�x�}߁��bw�Ƶ|�?�w?�?x��n���<�ü��#��!�DhPHdc��� eI�ߦ�p��|�|8ŝ
�,��o�y�.���7H�U\�Zu�(�Ӑ�d֧o16���)c�[#������fqila�����Z̜J�h�>������Xl����{j5�m]�!��Q:��k	,M�`�Q���(8���xG��!
1G� �U
g��[��0��P^�ku��z���aJ�e�@g��)��b`K��y6�=�!3��x��2Op3\�����	ҲF	fYJҰ�g�gI�Y�������ےX�;P����PШ|I�,Xc�x�T�Za?l��� (��ҰFi�1�65o�J�'pÐ@8����h
q�gxX�D�%�8Al�!Ӏ�٢����u��S��SPfABPo��m'%���I�dm�"��(�]p*��]	X6�3��@m@V�x	��b����
���b;�� ���$� �8�<Z��3PS�C�t1B���	��I����KaqwTR�M��ev�%v�<�򊏽X#53R;��1��@���(��r��M�F�M��J��[��T,7_�L��̌r�ó����CX.�I�h̋/=�S�<�`o��lj1�+��ߏ[� h����R&�<� �d��ٮ�R3��d<�?�aK����bM�{�d�Ь%�-1\�I��JR%����Y^\�3L��G���6YeQ�^����C:+ISf��/|��XRѶ,.�3�҈D��B�2p+����� �(c�"F�U�Pe��fP&h�!DF������SVE����@�,fe�&�\ylY'�{����ss�~.���w�����νoa�Ǹu�\;t/;��+GX?|���I�̐L6�3M=RtJż�"�	e��*'�*AF1�t���YD6\Ǯb<5��m�vFd{c����Q�#���("MI�1��	���`L�;���c��ȼ�g��#��яɆc����T��>��)�P7#˰�%l�9����T%tVF;)�>W�1�v�"�Y;qɎ�}�bP@m��X8�N=d��!{eh��#�n2��S��*-�F
���(&S�b1 WB���$�@�3�X��`~�������1<����4EM$/=q���4�Ȋ��,Pe��fI���hx��7�� RFQ�;�3*�Wg�g:���~�W~�����+���{�Yo���]��.�f�|�	eLYf�£T*������>,+�1�g�_�u�,Șo|�I�Ͻ�O_�đ�'�e���u�����x�/=���e����Z�H��$iQbJ�o���(,L�#�"�ҡn���$�.�Ȥ�h�d���`�R�,6�{����XL#�����z�����2Cg���<�M)윪#�]NQe�.�N�*��
UN�H)EL�FT���	�0��*㒢��6�2:�����b����oy��o����	^�&j>L�7�z�M�����)��E�ڦ����F	�`�D�)4HKQق܌��Ab&�D
��R�I'#��daQ)��p�LK�2��L�
2���g8�AkL���_T�f
׷���-�<�
C�i%*����!aw���*����M���xN���%n-���>������RDf:��3�����s��E���p���}�?��2�;���6��I˒�88ڶC�*QH��F�DE�O")�ē� $�Hc�&R�X��������5���6���7����Rנ�����;̶$�����K=�C�����m�˂r:a�V��
	���(��ЈBPK*tM0�GdR6=6��b�n� ������vˠ���ػ8v�$A^b��q㋏s��|7��E�J���p��oC�6Ƈ��O}ج*��>��wYz�骊+��2��*�m��� O^x���7�Ɨ��x0�_��4O9�c�}��Ge��*�aI�((��i1������Z$�1�Y K5f�rS,˦���&/#�sh��̉9F���R0������ܾ����&��c�Ħ�6�%Q��u0\24H�pP8�Bc�M�SǓ
S8v��j���$�u6�r{�0�7>J���Q��~��������t�.VOcu����,���Z��ZY�yh���#,?��=�Yx���+�-�>�Ͷ�.�5�~�̦����d�l�vٯ5�Co���&6L(bFLM�$5���� u�'����hڔV�̨�k ��B��E+ �� =R�`V$�B�>�j�T�FAD����f��͇|F6�9��ID�`Tk2nv��\_\���C>}��w�K����b�h$���B��|��/5j\��'��,6HZm�f��Q'q�!Y���J�}�O"*��c�c�g1sS����{GIr�w��{+w����9$ ���� ��u���_'�6�`c�E�&g%��J������Թ�r���Q�o��3g��陮��>���%�;~Ng��d�/��g��_���q���"�>��^��l��a05L�{�Դ
�e���ɔ�$de�A���}<C���適�V�LNL��ܠ>=['��>v]����[ٽ�B�Wؽ{7��c�<|?��::=�Φd}r�M�܄rD�)�z��N񃏼��w�������\�����߰4R����_D�ÆG���6�G�}ֽj�	�@��0��DB��q�<^���u(���c
K(lǠt�*ZiӰYo.�_Ö�����-G�_{/�܏��2_�4�>�#��G�ET=�m�(I��Hb�0��u���l:�M��e��f�h�-֝'�������WcOo�:<��H4SG�F6�S]HHh�|�����*�apBA#����fyv�sGN�����Z�����=B\#ŎM|C�`���Ja��Q�?Fa��	�6(��@X�����W7Y����j��'�%]��B�8ajl���:�n�4MR���J�G8T�t����0!�Y�v�p�Tf8�Dr6(�G�&)rV�T#	ɜ��t�c�%���ʦ��K�[-&lUu��1��e
��le��(UӠ��MC��.1��D���<��_����h�*ɼ�,�0��څW��"�zכq]�[�����W���?�?|�~K#X�6�;gq�Bi���f�n�K��!m��1�C�v��L�"U0i�]�&q�tC�ș3�����-ֹ��o)c����J���+��}�	��/��?�#{�z��h?�샨���'���GR�Aw��gq�[�ɱ'�'�"�i���f�����~�[n�+_���s�++�B��C
�*͖K^���F��H�3��n�LS�8ň�Cֻ�����i�Y]����e���d�����LՊ��yN>��-��<w���C���!-��k�RC d�� ��JB�IS���T%��M�k��"�&N��͛��n.���c��Cql�2�MhHBJR)H�Bi!B� T�V��B �Dh:Z�@y|�����`I��!9����j�X~n�ᰜJ���+oa�ʓ*�5�Z�!?T�A���e�r�RD�c�����/b�k_���"��#����ه�}7K�I���1������9���ѷ��f�ca�9=�F�ș@0��V��1Q�0L�ł�[b#�t�N���rc�QBT*��(��z�:̆1�2�MbzZȹ�l-Gl��*L^q%W���h�w�ى�p?b�^��ъ
ã�I�>�a��ˇ��^X� &�@yA��A�0���[y䑟�%��!�V�lv\����a�q
=P$�Dj:i��F1��cJ��3 �N>�H��ry>���)Ee����������qiNRk�Q�q�t�~��S�~�������o�ĳOR]_bch��7�Djj���@o�Ϟ��?�.xŝ�=�Wl�ٯ}/tFml�뮦Q�iw=������>@+$ҡ9P�U�v�aM }���G	�J0m!�w���F:Z�89��
��L��8�/0�.3\����^Fٛt68��wy��~��>��׾̘�`*�S��'d�߳D�$R�DI�@�*A�I���B�`�4�;^���^�y�ŘV	+��Z���tA, $F�1�Y�'1I�R�2Ҿ~��T�k�g�z���?s�e��xj�g�}>Sc���<�F�����
����ǋ6[T���:�cPo�8B#NR]'V:�DQ�dG*e���o���؋?����Ll�L����k���Sx*�n�(aњ]B�:�iBf�mR4��P�L��뇔j#�����L��&��3��}A`B��*.���#B�J(M���э��*���T��c�Z�}��:>D��0 ��%+��s�+�b�����#�����AA�P0 ��U�	�*t#���̕�x�;�K��6>���b��8�>ŮG?��,e
�#4�W�[�X�e�DJy��=�0AD	F9*��8��&���Uu����Ч�(�l�ȩ����F�Z˖F���r�c�i��-��/����p��1���"n������Xp�繿��3��M��RC]|�~�r����۶3y��=t������*�N�@��[�X�޹EF���KD1���Q���>�.Y�ڄ92A����%��hQ4btC",?��V�̬�V��O?���~����Gn��2�3�2�A+B���ef��*Pd��h�a݂��	6��.^��C�B��0-T���.��?fj�.B��	�R):��Vy�/�R6���o�|�K_���Շ��:|���ᖛo�^��I��ǎ��O�������x%GO�ة�T�
�����&Y6Jtӈ�e��zk��]D�X�*Q���9y���1�Ml�U�3�w/�tn�����P�!Q�L���5��6����bV�����^z�M���a�	V��?��<s�n'@Z6S[�XY_��M��y�b�\#e��A�Ld,������MC�Z�v|��g��MՋ,���jF�.�J�A2`h���>�vo����<z�����z�o|�o���`�s)�}�T�.���	)X&q�'	�f�BE�zi����?�m��y'�?w���#��骘N�G����΀���D�j��ɧg�')Kp� ���lR)�Н]�E[.���z���YL&vnfz�f���
y�T'g�IE@b��r�eS�w���W��ă<y�˸�o��t��.�0� 7�N�-�s���Ua�[��C�%Yn�+���檱Q�RrC�D��G���tܕN.�Q%����J9J�C�R�0�1KC�.��E�o��C�`��gj|�����D2݂J
�W�4�{h�1
[��"BM��V(졐4I��2MI�iDI����!t����
���5\�+o#.TA32�HA�$s�6}%��F�T�=��{�79��n�����GH\sݍ��_�%�fN1R�'���%�����B
ֺ=����W�����n���.��qP�T��]���L��hx���������V�J�L&���K�m|�ޯ�vb���� A� ��)"@�r�VC3)�[^�fr�8�n�b�N�+F�c�����EtGG�:�p���:�*0]'o
T!-���Y��2�̄^�@je��
����'	u
��>=�z�ǹ�s8��:*�N����fb!�R'?Z���~�ɿc�ģ��b6�&���S(Fre�a��x8���3�v=�5�#�Q8�4����v=�c�>R�ր��d��%�ÈM�J'��V��b��p�5p%�5*e�m� ���v��d��Xs���(R�ȧ �2P@$R,��!�ﯱ��G��k4-k��nG�$E?~���O)?�#����m���{a�ăBn�)�:�H��S�°L�  r]z�N�ĎM���=��ˡ����:I�H������f��gB��4�2\��1�Y �:����c!�Y�@�Ǚ��a��6���Nps����y�N3�`��4)��2	S�nڄq�@1��\���x��:i1��"c%QJ�o|�[���>�Żw�IHb�����❿����k��Vn��eb��y��~���������"�|���&IR�w��=��S���W_ž�{��/�����7��&�f��c��'b0r6�n�����=E��E>J�(]�1�4���Kxխ|�����~�^��_'"��[�^�Ŗ�q>��P+���sE~�mo����6��E_��=>���;���L�R�VG3(�E4�d��IB`�4��"v�n
E�P�^�M�%vm���'h��ٶgJ�{�IƷ��/��/��P(@�u%�.'����?�x�I����4�8@!2&Z��t��̘\��a����c�.MT�E��Ĥ� q"�E`�y��KN�ĐرO�TB�QTSE����L<a����M���ᷙ�1N�PV�P�qVzX	�KE�(AW)Q��@e�.�s}N��}��I+��7U�R�c�y�o����c��&�3�1+[�i���y�������4׾3_�}t����Jʞ;o�б�����:�\ęA���̈́JÔ�機��Z���2�菨��y>� |�!�0B7$Jyb�7h��bj�<�ء�Z=�6�A���2�r�مOc,�$�,� ��Z	3��(���\��wb�5���в�2�S���y����|��\�g_�W�� ���?��#c�����3O����=t�&"E�)���㖛ndz|������o�������o�����OR��pϵԆ�|��_�׾�����A�b��CȐ=A�/���kyky#��� ,��N��W��ts�.���g��u�$5�za@��@�1/<���
&I1�S��X]�5�'ݱ�S� =�����R��b"YĎaLڨ���`�@��t��')I�s.o2������S}��ae��r1&v=��y��9�>�����5���d*j�����ߋ��/��;���Id�kI��Ya��I��j`�:V�B��H2�I�@�Q�"%6F�)��5��@�0����~�>�g�\����!=����/�y���z��:plr9E���z��l0������ ���YOd9z8{/`�<�ѭ;��o���� ER@Fe�V�4�54A�T&V=��K�.���qf|��߸�#�W����_���ߏw������2|�eH�]q=���"s��O���]��fh�ʅ�������y�o@�@�e�5?���@�A��fyD��nDGȱ�C��4�7��;�h�ǵ�ŭ����E^�nJ���2/I^k�2�q��b�q�0���%���?��݁�M�᠑G���D(��X��He:)�V��~�c.��
���j~�p�Tc��o~�^�͞���|�ӟ���	����8	�7ژ�,�<�cZP.p���� ��ƬqSM7��
�CRQ�[�m9ڣޤMs�b�n#�M��	3�q
K���������������=�c�����=M�z��ƻ��!v��W�4O6r����J$��!���$:n�������eZ��.Zj�O���
R�b��P�6NYE�Z���G+T�D�-��L�JL�LT;&���^S�5H��H2�t��hqH<B�сT�if���,0�4s��A���*&)��%���'�	D�	z΢��)�=d��M�8�`�}'���$�>�������\��w�z���+^E<� 7Uڲ������?q�?��m���?q���}�Ar��o���⌌���1�FUB�:����胊 UhJ �H�"�>��!BE�@!�-�#P#�i#^��?��0���w������S��%��[��;`�4i��މ�t���=��|��;z���)���?e������}��H�1dXn��6_��苘+]�ig��(A��Y-0H;��Tl�����Q^��,�P�m`wW)6��k�c����9C��$Z�8j�,4W��d�%�4UHP�!%
�0��O�2A�(��ֹ��Kؾc'�i񒗼��g�bh'��?��3|���ݿ��|��@�YA���Ye}�뱱��s�=�/��n~���ݹ��MӬ6�(!0���49��Ρ�.�>��6|�]^��9VO�������Tȵ9�k�&�:�Tr�3ّ�s���9&�B�]&v�Hb�j�eSGKSRM�1��Q�&C�2����R�2c�8�C�E��n0`��$�������ns�F�A���2���)*ԫul�B�\�loO��$�|m�@"1L
�Գ}>�  �i6�ӵl(���t���"	 D G��e�l��"S(Y*��FG�����Ӝ��#��7�����/#�Rzz�^,�v��"3�����_A�̲����/�ǖw�6�NC2`�� ��0F�	q�!IbB�b�0ίc k.h}L�����HTJ??�F~3����c�q��X�ma���9{��X�׸ڋ9��A�v�U$�꤅B�[�BQ�Q/MP�jl���UlOY$�J�;m�'/gu�+Y~�o�|���ⷳz�+Xݴ����i���Td�g[���hZ��lL7@Oz�V�#tE�/�X
V�����Z�@��-]��Ǥ�"9oi�$	R������5�R
M�8y�$7�|3��a�&�^{-�O�FA��g��=g��j�1L#�AH��,�O�������3���[��?���_Iw�ɄY$��$�A+����XJ,EeV��Q�u��t$�9Xq��I����
ֱ���:�4���>w����9��2G�1w� ^8G'Z�Qpi�^�'Gq�/B|bbM�D�D%�F�$�Q��#�H�(����6:�:5�a8����J�k5
�<33����E3z�.J@���E�)��BCJ)@� đJ�E�R3���yZ*��(��\j���31��Vcze9��"�U6�*�Ģ��,�e��V����Dyi�ti���c�p�)id�=�R���H�	s]���>�ױ��c��e�� S�r�V�'M4��DM��4�U�g��g(4��Eq�D��M0���ֽ���V}*�[9�ܠ�G�m�Ы7��.��J�A�C�'��\����a��<��ؔN���V�A�Si�3��[�fe��J#yN�n!wͫ8:5�{/���
�hKk]�4}=o��`� ��E(b��%v�h�"�ۧi��t;����E�F ����ن���]�f�3B�����	����u}�Q��uv��I�Tbff����-�i��m۶q����׼�]�va�6�����ʫX�h�X]G�!DJo�#
T�R�����\~�<=� ���f���Ckv���0�ހr.��aT54]G�)Q��T�ptT���:v*H	E�4a1\ _�&�w��@s
O�(F[PE��Z t4n����CGY[l0�/�s2�B�Li�F?%"�(D��DIӀR���y1�J�J�L��Bh�8!ɡ&�b�4X[_B�B�D�2�Xe�+�4FI�&��P$B�nc�Rе�n&IJ
R]bX�m��.I#eL�[�U��V@$`i)�1��~5O_:t+�(������(�}�af�i�PܿTJ��Kq���0���}�!�]���;B�SEģ]��^�Ve�]��K�կ�9�SX�c�W]lNb� "J�҄T��}%��8O|�ԯ�v\�3T���Nq����h>�uXn@�ʵ�)�N��(y��i�*t{�z�4�l\h@!�s&�B��B M\�`�3�ň\��ghu�*�=�8�O�� H�����.̐M�x/`xM.6#v�f9gl����bje�5Sc֐lh)7�:�`ב�ML$��!�[�d�_~˱�R��)J)�P�i�X\\�4-,ˡ���Y��%l�fuu���Q8/�8w��7oFHI��,--��I��u��[6a����g?�?�_�U��5�LL����y���J��y����a�%��d���[�y/`ة!��L	���hcx!��"�Xh�g(r� H�z����r��n=��a���N�l�zt��#�p�ۣ��!r�n�N	���]�s����tta��.�|�v����P����EJ��P)$B�0;���0v�bh�D�Vgnv�B�����O�y���*W^v�bad^NR�(����7�~��:�$�����+�H4T�]&	�bj"s�W0��4���ӗ�U������U6=S�hm/���\��P��������>�,#^�w����x�����^��i�t��C�'��}�ox���g�C��I�6\�ŗN�ӯ~����.^��s��ހZ=O�K�>�]��'�z�6|���9�җ)��w�W*<ـ�?�?�f��T�y~c��J�u��9�xL�s�"�y�ǅ��rh���a(���ET�~^��9����P�s�]��SO��D	զ�e���[�T�+��O�kG�>��9�A�p�l��\���sk��G����+�/��l�l�yh��Uu(lc�/�:��|��eΟgV�G	�a��^�n�(cY&i�"�<�Y��hz"+�Eֳ"~Ʒ�0J3�-
]J��_>ǿ��0>6���4�<���a�n�ώ�1�a�~����?���q�1��.2�=���楸&$E�H�6�ɑa9�i2�Ð�W�̀^�������b�ݯ���/�>7Gί����i����6�����Eo��������>a,"��n��e&��9r�( ��giq��1R��nb��+��r6�Hc�r�B�X�^��R����_���������
�@'!������E�Ǟ�X�.�1�i�.O�LP"c��P������ܾ�vm��"�͜ô8���GaJ��3mO3�L&/u}V�
ֻԇ�i�.d��a�>��@JlS�{RL��4*A��qק41JWx�
�{�8[�E
���S$�H�+<9����	�z	���'	��F{��23��F�2;Ӥ3���h��z� ﰮ���4v�m�w�l���($6��0c�,W�"�9�����P��2��Bէ�5q��T;0���@��n��4�mAM�\�#����vR����δ���!�����-��)��<�R���C��(M�p\�r��15����ha���s�k_�ںMf���G��d�����އ����7�?��Ǐ333��|>���$qL����S��=F��?})%�>�,�{�h��`����r���1�fOq�2��=5���9.NtvzkXgNc����k#��=rk�Vϑo.b�/b�樵��76���g����1v��w8����'ދ��OI�?J�;=N�4��g�r�a�����5�@���:X�C�\B�l���=���q�.N�&M��ޠh9t�]T�)�*�*�^�b�t^��{C�e��j�޹�j��8�F�}1��G����>��PA	��D��d�M�<#$k�M<��z�?z�͙uB� ��)���L
�!�ހA�ş��$4ٵ1d��Aa�
Q���B�as�F�e��
LZ)�z�()�9EE/ T��^�mE�EA���3��%������G�������W0<<Lij����~�C��H`�$.�Mr���bh�w�|{-�֓94ʱ`��P�Ry��$^�B��ѫ
��eV��(<�He�\�J�q��:r6a�7JE�T�E�3UX�$T)�ṵF.1���Q���e��/1��~�J���*�X���H#�9�h��i�ǈ��./��}�bj����칄�W���Pֳ��7�R��@�uM���ߢ6T窫� Ib|�G�3�<ý���\�?�A�n����4J):ć?�Qʥ2���9q�8�^v)�i ����<�У�ܳ���1Μ=KG(ͦ�/��6Y�,p�ދX�=GQJ�r�\��q�̟#�2�P�{8^�)�D`D`pCT�c%`�c���w�����;��g�6�b}��y�U��_E���*XZoc.��#-���RfD�R$���hvI҈���"��K}�����M�m�J�F�h����	☼mG1�vύc0���(�v�X,��RC(���{�0��c�SG��!����g�~��������6]Σ�=�WP��bw=b! P\h���nbw#ȳh(����"�%(��+��:}�����9Ӣd�&ӾF9��m�S��$c��Dl3�$��b�t���]������n�૟��G�dוW Ky�N����q�=���I�@j����1R�f�q�%=�����ƪ�X=s��ӏ����0��/������Or���w>��S?�M:D�#�t�M;�d ��L"WIB�|hAb�&�����7\�T��in�@A�!u�acn�#GNf����:2��c��n� ��R�MB�Feǥh��i�2#ͧ�σ3Mi��EO>�$�\�ӧfH���b�C���|�?��?�+����8���DQ�`0�;_����q����_��_���qz�t��aH�T�e4M'Jcr�<�n�v���Lo�����B�M�WjDe���O1R�Q�%�m{rQ.@�`&=CHl�B�W��T�H5ttL][��y7�����"g�u���[��7��~�P@/�;)��chs�<z}���!�j��;}� �P.�h�x=r�M�R�R�fC�$ #?�V��m�nR4&�Bu^����i��DI��2LDI������&(D�'&#d_��R�k�4,�y�@����]�b����r��Bz(�Cj)F�����hF�*�Zͯ38q�����ì�p����A�����Kx�rF�O<�F`+!L��N!H��:AO@/ґ.�O=���#�*T�"�T������$9��F���lR)�7S�4�E����N<���O��o�C�����c0���<� ���_���79q�(v�L�YPĹ ,@ӿ.�JQ�s��ʎ?�%-|�'4�b��uRS� Z��z���
�R,����/�
��`ԫt���:��-,Op��6�<��T����V)�a�i��?�'���Q
8�eY�a���:###�E|�gdd����RJ�nن�eG{�R��{��}��a�:��!4A.��왳�p� �|��)�0����I�zč6�C�Ȃ�\Ц5����qh��LI�15D�i���'T
� �S�(@j�4HR�"!�-8��?�i.z�Q�/1rǭ�W]�9�&���	���ˡ�
Ķ$�r�I!VT+5� b��.ab���S)���gtt�ng���K��H�AN�V�^���Ç�� �ʠ?�I����r�B���'���'���'��P�D	�ʂ4!�t�e3I�Y�@�)fNaZ'��P�D�.JF l<���Do m�	;G��#��H�`��1�=� '��eV���_�/ֿ�U6��{G�>K���.�hg���HF�~6}�(0�����n���(�� l�0��폦!#!�����`��|�Q=�R+�7
�o��%9��%�8�OS�\grz�w�l�&��/��� G��EV��]>� ��� ��Y�N�X&���]���%"/M(PJC��7��&��8&����`���̇(�g�;�V6��K:��\N��o����Q��F��7p������Bf�	B�,h�@�l��j����a��m�얛��7�EE��ɖ-[x���q]˲X^^fnn)%�\�������_���~�{!(�sHMf��$A�ׄj�zݝ�*%��I܄������q�0�/���`�-W1�G@�O���{? ��:w�B�-�Hz�><�B
#P�JA��1��*"�t����W�E{����x��lgx�49=E�u+ڔ͔�mF���GObZ�<��Zv�Eq��NK7�|���yVVV(sl�4���)�r(��+���4tt�@7M�T�T�%�j�R��ne~��z��k�Aq���R�g� �*�ޭd�묩��A�i�$� aP�I�<�7Dq�A~��5�;m����#����6l��!�0�o|����`=��p`���N�c?f��{x�x���#4�L��6� *��3�"~Zn��!;JyZdBc ny�n��#�}�������V��g�P}�-D�`��dKc4����T�)�%z�Q��G����w�f��������2:Ǝj��et�������!�'�_�����)�-G,s�Q!M�c�$a]B��.�.��\�e�b`�=�dP���h��-����#4�};S׾������r�w]�(Im�R)�R�`��Ú��h��8~]׹�Ɨ���z�kx׻�E.��Z�255�=��������֭[ٿ?Ap��	�쿈���ZCGj��Z����/��Ǟ$U:�v���uۦ[�m�O�|����l�`���f����魌��EԷmf|���\�����p�g1���Ҹ)e�5x�̵|V~�8�o�����B��IZ��q���,?�#�O�E�%���j�'4-�z�$�UL0���������2Az��g�� I�����H$�c�&����u�r����"�b���LL�bX4�f;M��c'Y�������2[+	���$�³���i�ιMW��~K�2x=B�:�%h�`	���Rȳ���Pn����.�=�=�՚��h�%��=��eT)���l0�̆��q�I����͔���>�vjP�$[�ɞ�aҮ�[��,r��S����&���XA
�ДN�$���%	h1H��B�"'ذr��;�Ɖc��㶗���v�3^���w���{�]��Q��u�n?��r;��ͷq��[�N'��|w�S* �ub	�Yx
b�r��xn��lC�)�M�	�*ď^?f�����YN��;]�C�
a��4����??z���.�̯7��������G>��<��O��+ ���N��y�}�K_ʟ�ɟp�]w��O~���!�(B�4���/r˭�b;�����E�ydE�.����0$G���X.��\df�n� �{b]14>ʣO��E/�}�a�<��.iUk$�8� ��L E SГ�@(@Mm��w���0��e,�4��t��=�������*�(��n#�<��2�������_(��v�E�١P.R���4=�m���Yyz�����s
����fNG��F�������0Ke�\.c	)a�	y�9A,��6NSӗ:�i�*��*����0p{&6AᨔS�Klڴ�V����:'fO���0�7�5Qf�Ra��I.�d��p1�]4����ʭcLL�@>�����S�S�$A�FM"2��@�Y�,M�(�$��T6	�.$Af��**Eh�0���$�(D�����:�q��,�t�<��ny9����檋��p�4[&zGY8�.�3���7�r=������@����$a�$D���^f2j�ĭ&�!���~�
$�j��A"REy�;FX�����ۙU����"����m��F�<F�r��+�k�0{�?�؝�.�dii�������"M�0M^u��9r��`�����}�0i�Z��uL3�AGGG9v��&��7����y�̲X���d�����il4q�t3U�7p�{T���ش	a����[���~���>ő2z�����KU��T��T������rD�vQ����]������=�y�{����Jv�pW��5��M�0?3G���4t:�b��s�}�(Li�q����e�b�;���ƙ�g�Hex��e[�O�X�0`ue��'�Jc
��R��i�i&j����M`H�i���iyB��9 �R$d��X���J�$�QN�!�
�XQՄ�
�������c;Ɖ������w�'N�h5�t�i'��Q�-3�_`�\���F�x�f�����-�*�'��qr��%	S��2yZ"@3�����~@�f0�P	ife�:	�8�QJ���Ć"%�d�/�����Y���׾�-�E��cs����o�կy���&Z�~���o�#�{/�f�(0��x��4]'I�"[F3l��+����f�@��N�h��BC$Ui��>A)��t�[��ʈ�����FF'��k%,��>��z��"@�*���T6���r8p��q�$F��}�/��k�EA,,,��O��3�P��%�"��� ����WTk5^���CӲ�<�=� �4]G:%li�]��F�P ��
��g�.7�fHN�pb�/��v�䤉H��D�6p��P����I;r��y��od��[�]5�M0Q�t����P��.�(*$���r�^`"U]�A�0�e����a[6�nò�Նطw�irv�$��˔
9�'����]�Ӳ9z�'�a���R�a$Q�La��W�(��E�"N?;b��R��O��X�l)�ۅ��b��d�$,�A�����p���3V��s�E�xӫn!�5x�^� ez�H��qp���}FF�LJ0\���=|9 �4!HJ��B A�1���%
S��
l�-;��g�!%�۶`�;kR�(E�I�@� ~�7�461�/rH��+_�
����&��C�ڶ�k_�R�'����+x�Ǐ��.��(7��
^��_8�AI��.HI�t��b�uҊ���N�8A��Ѭ�(N�6ȭ�K-"�D#X�!0XY�����<��O���~�W�����,�[$I*MPi��#"dZ����⋑�DRJl���/$MS��:��r7�t/zы���Kq�癱X,�ڻ��]�z/��ѴL�~�1�B�B����}j�n!�I�x}�8�1���]np�����_�P�\�����'p�M�+M,[Ȕ�3(B�nAT%rT�HZT�����<��_����.��0k���,~�����ظ���OS�=R-�*c���|?)d���Jy����aQz�.�p��Y�R��kU4Ӡ�m��1���Ur9�ёI2?7�̙�$IBe��L)qE�(��e��D*��D�"��(=_�
A*2c)�Ehaʅ"�>�S$�=�w�1,o4���Q�:$�z	V|(�@����Lq��aB"
f���	�7�g͘��~	�vL1\����S*A� 疈֗0$�D�z�F0�Z�X�Ј� q~OK�,� $��0�4E$qv��f�aRtb�$%$�m軔�Ð�P����5�������b��er��Y
eɉS'���>�#�����<���ׁЄ4��jI�ىX��?C��)Z�N�13�����3�������S�$%r����@�W&*���z�1����q���y��q���N�? N�S6MҌ�3���v���%��nv�II�$<�#�"z�qc�6Q�$	�^�T)�8�u]<��9MP�u
˱�=����(��kĆ�3�6*�n�K�K��E�A�=�0㎞�9I��`e��U�
xJ��7R�5Y�1Q��i��p�v^r��Q�{���8J��L���}� ju�z�c�,S*٘�`e�B�t��7Yk�S2M*�
��cc#���c�6�c㝷���0l�K/����w24TG�:�&1t�V�E�^�V��j�0�RC7��>M����5A���^& P�=+5��g��l�9����,@E��"�a�����P�O���s��4q��k��5"th��\59Ɩ�
۶�1�y��^�:_�^���_}�M�#<���$�&o��v.ص#�G���]#��8�7J�)%�v��
?�V3J��FA��ɠ1���Ұ3
����=�&Ag[
�y+��Ƕ���e
�GN��P������T��Հ?�5NΜ���c�z����7򮷿�v_H�@�g���N�s���m<B������u�y��e4zJ7'��XK	T@�ns,m��H\��Ra|vO��G�����w���T�o4Y.�Ϝ`��$�2'�0���q>@�$���O��Oy����'>��C�H��08~�8?�я��~�=����������c�&G�����_�*�����g�_����g���ФN�����'c�R�0M�ml0e�4��q��j�����ƹ�#�� \#�����>�s��D�Z�����(��xܗ�4�Dޣ�/�X��7WyȂ��}�GÔ��dє�s�VDXH)�G��F��ƹ�9�WW8s�^��"I0S�~�3��,-,��
��x8y�4���������C���J�$��B��$�,]GC�!���YI���])�B��(� 
�HL�6:�T0�w0,��R�H��T*U�m�֛Pp��+�M�uU�3�`�����̞]�#�{?�x���s��h�[FZN���|)���@�F����T�HiJF��)�aB��~>:_�G�G�(��輄ʰ��%I�e�e�X9�����U��c��b�������Ĳ���?���u/��c�V0J�S�g�0>�V̳�[���3x��1>�>>�J�F�#c�4�$��Hq&F#��<��T���$�&p�����A�� o۲������H���BD$q�P��ZN���j�7�ͻ��n��.���������/���o���o��;g�}�m۶!�`��ݼ�Mo�o}��ۿ���"�ӛ�u�T��F#4�b����M$2"&�*�I����2;�u�F�pd���</|���{�i.<�����e����\j��@�<b4�jqc�KX*mgiϕ/���u/#��fԞkh�p�+ތx�M��(ﺎ��m˅��ij�8M�ᆂ���Q�����Q�g$�Z�B)_FJ�e�l��h4��ju�l��`0 LR�V7�F���u]��"�ccx^��ٳ��I��r�BjI�]#����0��4��9Y��t�*�r��%dtiY��� 4��z~iu'+��D��0���Щ0�یp�!J�Ar
)"�<�W��!��.�w7�t	���N>�������l��{��M<��3� �i�NlbHz
Tb ��.��8C���$���yRI�%3��4�IR���$�7�ilt�b��(��F�m��Z%o�<�,G����?�qZ���ۯ���)��C�N���Ϸ�c�y��M`�X!L�vU�<���_��`î�عJ&eW��R���	^c��O�p���}�K$SRC�N�����'�>�y���ǘ��!�уTg�X8|�n��f+�A�&�8�9r�(7�t3�r�$Nغu+q377���a�a<�䓼������8###�i�i�X����g���|�x�+��k2�Ej�Q����maJ�#Ǐ�1��*�Y��'��3^*0tY�i6Z�I��	���?e�_����'����Y� n F�y�G�υoxk�Ό��ɥ�<ל秳G9�x�]7\��{�뮤?5A��K�w��v��E�T��D'uu6\� Jpr#C�h�FG�i�4,��s=6668u�� �^�#��ĵr	�i�[mN�<N�$�L��|b�(U*�(���	"�l���a�a�f�gR�yb��4t������OvS�"c!��0j�P���oA��v��	ZS�硚�0Z���'��F��/����gy��?��?�EZɯ��6���^|�Ŭ�\�;N'J�e7�\�D�$q�WIo��؏AJF���?���y�罐���R��u�(�&}(p}�����a��846(�e��E�]����w���F��.���M�)qӍ�rv�Gg�R��ÇCZy&r���Lday4� L�4Py'�0[&��n����Xé�bd�HT�Y) �Få�)��S�T��FE�S]w�/,���aK�b=���2�v�n��/""��'�A��O?C�Z�R���ؖM��RX�ŷ��m���w����l۶��%�����yv���[����.,�"�"�02hfey����߶�b�B������P/�H��x�F�36:�p�G~i��3�L-�3ur��S���ȹ>Ų��)�4A���?|��$6\r����_�_x1w����X[�_>�I�+�Gx�o�o����_���⪗��8�2�ǐ 4L���������ϱ��H��1h��A��E��@0<6���2��G�*��6f.�H`db����255����q��$�j�B��i@JG�e����FM��]�3��39M ����]'�S�z�Z5Sc�}'���fC���F�?h�sK����/e�X���!����]V�Vx��<_����?�ݞO��cf�,�4a���Q�X��0u�Bٽ��'1�`X���g_�3��ٶ�N�(4�A�ez��G���w�� 
��y�M����.j��M�p��üᶋ�����]��k.܃�����o���Y���a��VX�R�'��(sVO�z!�)T�^Si�
)�$E�PR
���/�H{�=bw��`u���~�M1����+/s<���e��c��j�'x��!V�VY^^�s]R%������y|����A��{躎R��~�W��U|��_axx� �ᖦ���ƅ�\��C^�;�,�4�zU��0t����e��#uေ�a���JEvo�Dt�h�r��F_)�#A�BߥHB�����$��:��MS�x�s�'���+n��_奷��k^�&���dUٹ�,Y�׋ٶg�$���9�6�~��Y=6�6=�C'm�b����}�NjCu
�23�7 �(����.+���*5|��Ѳ�^9���t�x�)�.�w���������Mѕ"����<��Gq�����r�$U�IJǄaL��0������ʴ��}f�\ˣ��ꃣ3p����q�~	tB�Z��k��?�������}2=|1��],n���:������E���0rì�lX1�MoC�M�t ZrJӱ��<oH�>YY��8s���@B�Ě�eU!Φ\��Ax(i���V�������N��Вˇ��w��y���e�����v������{>���ϯ�ڗ]�x%a��n���1E��6q^��K<����Ő�!2�C*	���0�|}_&�A@ky����h�#��
�"�#v�\Ec�Y��pv���f���)�s6�kǘ�����'Yi�h�[t�MLK�s��:���4�M�y�Y�F��4��?�����n݁����o�K�K�I��C���x�o?�яy����L$�ID)oc&1[��~� ���U�ǥ;�YE����ԹU� ������غNz�䍮a�:��M�vH��q�q��Pn��a�/WI5+N o��z���d4W $��ø���I�]��"�9�V	�;��;K�� �'�)~#@&�V��j7H��X�7��;Jrdi�^��g*F��(O�ӣ�p��4��hT�5��u��:���#o��ѸI!NP��c	tbR �$��lt��	�A���0a�<Kd�Gе�(A�X70H�|P�ocW9����K�@�o<��w�_������r57���Ӟ�>v5o�����>A׃�%.|����E)��5����26WǤ�C�c��YC	3�`E������!b��.ǎ��Nb��<sj��I�ќQ@"|D4�0,����*tC�]n���pٵW3�0���S��u���*"���-�X��Ġc��y6�1���Rb|�vR�����Ht��2sQǂ4b�����v8��]��3����y����8�1�#��
6�j�4�Zgz��$O��և8f
fO,`;9*�
��	|�4�_?�Y��2��������_~�/s�uב�)K�9|��{������{��ﾛr��;������ηF�����[nf�V�NK>����0�
�2�F�͛&��[Ʒ����J#>�S�3l\�kQm��ř]�T)m�Tb*Ah��vC6�y���E��at���;���,gd���9}�q��=��ģ<��cy�a���78���93�51ƌ�Q�א��z}
�;7M�,d��tLr�"�P*�,�]��l�@�)`�iQ���u��CQ�,/�a�s�+l�2��'��ӏp��'X;~��?�O��7V�:=�H�#�}��Ob�y�X,����T��̱a�h��W�n��5�
z��Q�&k 5�F���@b���j@��ì��<�k�4�����{����d�+.����a�}�k4V���{�S�����	��l��e�U�.%��8a��<5#fS���E���8�o|�^ZO����"��P��}�}���t[}��$����[f��Q���G�qH�>i'a�2�=����eP	W�����/ui�&ã����<����l�7Ήu�χfx�k�#.:ͱ�ÄV���|p�l{I
���Lh�+O�&�L�{-�s��D&�n�7��f��F�n�E��Nad���Go8+��M��7o��'  ��$M��$)�7o����k_�������[nᵯ}-�����'x���O�gO��o>��LNN���R��ͣ|��������^�+n�ǴPIB�|����9����ٶyA��;w�"t��ȹ�,./R��`8Mٶ�D}��d
���]IhR�
A�z����v�=�����'y���^`���`D3�����y.��Z'fО��^uѧF`d��aR3GѲ)(A�ߡ�w	�J�H�HE�&S����8*�j0���`)E9N�lW�ݐ0�qT'�G��*H��y��.�a0{��(W�>���� \���/�	q����"��������ZF�u��Ja��]l�bVk���J�lm�yTb���2*�A���ټu�R�g~p��Xfa�w}V�Υ�7a�y������3y���4ش�-�\�r/��6�8E%	f�Ș#�5���xq�������>��Sg��UwB���g�/�����x1f}�/=q�w��Eǲ��3.�X��A97��,�9
�`��l�BΠ�o���!o��71ӎx��
S#��CL'�Rۡ¹�Y���A,�M%$�.��S~�;�'zI���,����9T�%6�z�B���nc����Hm�0;�Tg�Ze�o/��l�����j���)���r6o�L!gc[:�w���9h�Ĳ-�� �q�qW��G�$�|EJ�8���v�4N�*�4�?�[Q���w��<�,Z��X�f��(o�+s��#�z�{�1[�'��5v�}^77���E
�2I��!@I�Jt"ұ:O�ʖ�&����F=�^�A���9T�ӏS�&
�mf���PH4��F�dm�Js���)� %S��LA�b�ɘ�IHK�X�d�P�4�*A7�l�A�r6�8����az�erJ�ǧ ��&�t�e�J�xk�*��Y���Tq�4tߣ<���ȥlb2�7_bF/�|����ѻ�9���	q��I�X$F�UfI̥;�	�h1�Ҙ��F���=���<
���jA=��D:ǫ�L���f���9:�������,%�D23{�]y�Hd��� Y��|�;Gh���u���<��_b�?������/���?y��?	����rr�nql�ə ϔ�R�-�A���!l4M����m۷S��$5-���C��Ѫ�l�}\�O�#V:�k��bJf���MG�|��l�ig~�*�"��p�b�S�\t�l���%�y�v=B�Lj�:���ٍ9�*��u^�n[,��XKq�r|���0g�A���l�*4�ƴT�X]]A�u�8�T�����?�)�� 2���-�(�IU��A�T��%q�����7�����P}�mcL���ivi�V�On�'��8\�R)����B�G��Ɖb�L�L"�&��3�*�̻>=�D����.e�5W��׳���س7{�o���۹l�6vm�ɮ��`�����j���o��^�=w�	?�{������t���E��H�E.i�
�V�w=.
"v1�A���U��sl��Z�\�|��x	�J��VNa�Zg��"C�ɭ[�;M^��B��:�vN��M6�0�T�tm+���mV�C���"#�%F�VdҔֆv�O_��U����i��� �2\qz�D�<r��*�U�b�VVػs���bN���Nom�g����<�/��W9��r��N.�S�Yt�>T$�t�m�$FY�9�t5�)~�ҝ;�/��b�s��).y�k�RG���} �F���.���er`v�YYa$�Q�����R�G�0t���tL��7�ҐJ�aj��TF�۲����s�R����M���5�~���-� �Vg���u��ZDfV�Jd̈́�`���f�P�nPM�=�4b(��)����ҧ�|���(����|��g�u�|�$�0G�9�F��9�m��\�F�#�rN>c�4:����&Q�� R�Da�Q�<�<� �/�&iL�5��3�(z��f���C�w�l���%�w��h��������0��`dj���K��!;�J�v�pM s��I˂s��ӷ�T%3�<��#����~�C��o��O���0���}�)f�?���{�G������[���6�,�V��+����0���gd�a�G�Ӡ�w(NL�e�6.<��Sq��*������K=�S�b�T�26ʥ7^���D���Z��Slb��I�3g�)����ك��=�&9s�S_�&k/<���O1���=� z�ǌ2�:�YY��6<�F����.�{�P9��쾊#ta�4IJF*96UKll�"�%�}�8�*���#���l�|'kZ��={T�غ�b�9�@�<��m<7fbh�A��p�D�v��@��F�El�vt��:h��J�G�$oz٥O=���y.��P����{?�%Sk]zE;WG9'Z��,܊�*��Jg�H?����DS�2�ΛȜC���� td�'�b��slE-W��
�
~���i����n��"%3����A�J$��1%���	�Q����[0�6�^�X��/B����LO`�JDSF����]��u
�j>h6� f����8�A�T@��^ϥ���J� M
��y��������>��'�#��6k�������]�d~�{6mgke�ٙS�nl0�m�����2�vlò�h}+�#�7�D�w:�����1� �@S����d3���,�s1��j��P�C�x1Cg(�\��>� BLW�Xg�(�(�8K}��OW�nt�}]��v�=p1]&�!�ހq�O��òm�T�8{�t�q�x����H0�Hz����O5�$� �4td�D��0���ǀ���~�}#cw����Ss�Ԋ:[�'��..2�s��]r^���1�"7@�h�j�������Y	˵=������E�DY��D���8dl�Fxf����[#�JVc�,2�O�[��_k�_]�T�P�F���2E*��1%3O���`�E<!YGb'&a ���ʳ�l0U��� /Lh�;��W��{�QN�9�ů}=�hx�>�H��.�q���#K-θ9F�K�N�|�qV���;x����x���cpr���z�����Ҟ=���2����/�zn�եu��X[���0O����s���l۾�fǧ���^,d�yV�!D�R�.h�>;kTwl�}�����]��uF��J�S=�����q��:��2��2"J�R�\a|z�f���z�\ċcZ�u��!
p��D��Ѡ�n�������ngT�n�G�����z.�f�sgg��=:�>�+�����2�#�,�����F�)�����z���)�./��~ʥ�/AJ�^�A�r�PI��o3�뒏b�T���J%C�$Z�*;�|\3��r	�= ��1+&"�Zk`��\r~�OQ.h\�V�T��&.���*�� ���c�tg�%=��p��lr\��6Ta�eb��I��$�#l�a$]
�G�X�d�0C��*��e�΀Z.GA�(�7�	�;���ڦ*%F-��Z�5jf'����X���LK4 4$k2b1籘�C0~�x���I"t��f��P�Wl�+�Bʄ�j�R�G'�u�!��p�$q���)MV)Oװ�윁cJL�����-�����?@�r�X	[��aLϏ��� >��{_u'*_B�]W)BΜX��O]�RT��=��w��|���Ux�y0
�EY=e���l�*LPh���##�
�e�W�ٌ��끊����K���kXo�8{�,�N6�NHC���ʔ	6u�y�������H��S�N��`�6#z�FI��m#�� Jۊ��t����lێ�i�%��;�F����Op��GY�vp�LN�1�e+��1�'�0\+`�$��L�8��D
�҄$����t�U��G(�(-[}�����3�X^��1�V�8�����=���s�U{��i6Z�^�B��LO��Wx]s�K�2�q�HDJhJ�Dg ��
�/����y�4��T.��V�)MC�4lb\�5�l���0�I�8oNa	4�ʛx�G�g� }P{�p�R��5�R�WG�D)�.�-�zM7P*$M=D? ���ABO�R"�?z�Z���)�&^f��I�)����^!�L=���q� ��g&Rh��3���R������wq�ܔ@���:���tr��S,�`��� gB����� �soY�ߍb�b@P�1��t6ֱ�$h6�|���#�'������-cWNU���-���o��[������SO��O�td����G	ͦ˩�K8�����7���D%Oc���L��g�w���W;���f���E��*d�+2"���cd�w��}{�;�vBfA�̙A�������O(]�R�Xsk�͢Aǈ0�yd'a>l��YD99FJCD!��?��En��G8Bc��2�Z�X�
�\}������c�?�4��;}��'���P9uuuj�[��
 $� $���q��`��	N�����0��1��ǘ`��c�rV�Թ����r�zr8y�N�;�>ժ��jU�}������]h������J�v�c�ڢ^m�iw�RE��J��4ݰI9Y2��ja�)z�	����
��+L��ĥ��<��T���n��g�23�̱�`(]TŠ�h��m����~:�˭""�����ɱv+�����≐ o�ຄF��\Y���(2IT������	S"�2�0h���8qd�6n�@�*��j�4aO/�t��!a�ڣN\C��c��u}���]w��𝯡��{������.v�y��@�-0W_an��A(e��B���\ˊ��X)����M4��F�!2�����v�[=d!|-MEd�T�T��ڿ�Jl���/b�����j��G����෠6�m�K���7������l�P��6qr���7��a�M����� �7`ceuu�J@��]��lq]��lk��~Hsa�_�� ��g8=9ɡ7܏���+�𘹺��D=va��_���3�E=�TL� [5XnVqL_�����'O�ac��[�d�`�"�DH�b�Z
�evl�0Ӵ��ŕdlL#'F~�8#���@�c��p�O3�^�]�e���e�>{H�}6b�l2�����}��^�i�K;��˛��͈��a� j�A� _�� gA�i�����z{��rYl��P!��$�.C���(���qZn����>Q�%��,-Σ�mZD,T�9��Jƴ��ǣG6Y_w1Je��*�n��7L�n�9zO?Go���J�DDt�a�QS\���Y��9��8�[�i�,I�ompX7��T|�#Jq�R3F��q˂�&��ehI���L�����AߏI9)�R��D?��gd��t�b&�E�%}-��N
S��֠*�n�n����,=|��S�io��Wb�Y�K]����B��4ф�ņfs��E���*52nE��2J���z��9��I]gjǛY?x?�� 7�61(������88@+P�y�%�w�'�"�n���V���t�^����$zz����im����z,�5�6Q���f���G�������}��x�	~��9���?򑏃`�&y����A[蜜���U�Zk����.�c3�H�J�tFRK���b4�CѴH��(���:�|�L*C1�P̩8�B9�e����~��rD�h�"I����D��%Mqrf�Q�A%�p�D7EM��3�Wfo�F��@i����l� ��7h�1ž;
Eʫu��(}y�b��ve~15�h�a`�(�y�%�� t�|���Hw^ k�nϯ�l�D� k#@�_E,�#*5�F�#\��ԛt+hJDD��Msjs��ϞB'���@o#pJT�?j�Va�L3'"z{,��������B�OM�����uD&C��Ah�����Q'=���2)uz�E�F+�X��1~�V0"�~-.��qo�����Z]��0?���e��
�8&�_b߱�������;ٱs;�=�dR�i ��l�N������d��X�&��Pa���L���˜\ZcYwW�Ĳ.X!K"�혬#�N�(2�jT�<7�=&��@�[4"I��Q���uQOD[CK�J�b-�:d�i��e`�8#�􌎠��l�qk8Mi ���!�v1�k�t�;�����`��p��h�f��ѿk'�;���``�:�K3�"M�~Se�4h�>�sO��=C3�\���5�=��Q�����@�Vy��E&��i�g6	�kA�;�Zq�՛8x��R�ӈ�c%l"�*qm����@lJdZP��mCq��&iO!�!�t�a�8�BI�41�ׂ��B(�#S�b�c~���G��>q�K�� UΡ&n����0:!"��q��
��i�r�T������(sK�-��^#��R����Hm�J)�J����׭�h,�##I��hA��ȰK��†�%cLh�N+��np��$W��=>Fo_	A�PTL�!���,M5�X��Ã��v���U�,3�m��ё�AdD)϶�sk"]0ZLn6Qb�T_/eO#�4i(4k.�n��	��e�F��C.Mo�[�P��Y�~���>�m����5����r�֛�9�������%|��	{6��yk�BJ��s��@h*�P��7��������#�4jA����q]4�Ə:T��v�R}��2L�����k���,3M�������Swt�&�P�� ��h��3�0$�n�uT�Q���l��U7q}����.B	P���l��?�(�zHiiR�"��Z:���!�᫂��F�cR�Z�
��/���Ҿr�+W��� 
E�?���>.�� H@��z��g��=���xnr��P'�Zd}n�!C��uڑB63L��X�ΰ:s����|�Q*_�:3���<���^p�2&ah�ֳ�l�e@��1M�IZ�&h:��+*J#�����$)�-;��ܘ�n�M>���)��#e2�z��j7@z�D�Z%j�I��.(fK��!�z�]��n����PWuV�6�w�X�J�J����\�j�X���ؠ���Bs�Zs�����:W��pu���dji���e�,5*,.��y� M�o�i�&�N�F��C�I�L�"��fciuq�V��Z��J7b���Xn�v<.K�6��S	$�E�)���&��6����V]'#2Usy��������]�VLe����6��dY��拼�y��72�};�B!@�ԟ#X�R�@��g�UU�Zj%���-����6;;ͅ��y��e��ݼt�n�M�ql�n���	,�DC'_�QnV1=EI�ߴiZ&�R�i�Y�;�R~���&��iDĺ��r� ��t�j�M1�ƈ�tW(�-��{I�9=KڱQD@���l. �*a�S���E�U��,yo��it�%�J2����ؓO1�����n��{�<o�� ݫ�p�4���&d���A�V�8yy���z:�9�"=��+�>���ⲦnC�]�'�e������`z��؄�%�_F.�Ҟ_������j
L�b8��I(A�L��O���L&�D�e�Bp��vΤ�DȨ_e�$ٯ5��.q&�d����
D�KE�G7��Uvf��mT��\N�H5@�hB�d�f6\G�|�X�����J�]g��n���X��LJ�9r����N����C�.�Wb0��'Ջ���d���`�T��Λ���q��r����QL116 �0�˓W��)
��y$9!.�t�I4?M����0�gMh[�N�����Ҍ$�`T�K(b� B+���i��F�C�'�%f#D��pc�M#M��A����Z�|o~��������P5=�ɠ�֮)c;X�|1�����p�-*@�������h��7��-�W+�t�-\��<�ԓ,--��uL� �cbU��i���71� -��~���Z&}�0�Ŭ�&K{^�ty(	�Kl��-���N� ]�\(c;>~��0�i��T�\a�V.���٧Y|��t�͗��v�,�f���,�>�>���7q�>ylZjUS�ZL�
�
%Ӣk��v�,o�i?��9.M^����br�6���]�'h�6'g֙,�IV�Q#A[q}�.�O����>+S��PR)�l�3���2��FXtY��3:�G����
2��A'���`h��ҍ��R��Tpv�1�+W8�#�`{	��q��a�,z���VpJ=�2c�2�Z�Ҧ�[B/��-�J�Lӈbz���1S��}�����T�F�r��P�Foe���&c�*��u��URJ���rTt���Dc����^�	����Z�ǩ�(7��7jl�i4s~�����e6�(�.P�X�ou���e�*���/��Qage�n�
6�{)+)�+)�-+�+�n|���A�����uRMAx��0e��K�R��I�
TK%�]�b��j~jH�/���<�7q��k�g3H��n��t)��I��脢r��Ο�dhh]S��K�.���3<<�m۸��g?�Yr��qL<��G(�|�q��#��{8{�4W��b�Ҩ����Ĩd�5r�u�n�N�m P2i
��8��F]dY�+�!Pth*B!r0L��$�gj��3 "UĮ�@� h,r���i>�8��J2��dA�-r��f��)�k�4g��-����D�GU���DN��b*�,d�T�::�N���Ҝ=����� "_�g�3�("�c<��Db���A��ƚ�,�I��\}�4�|�0Z��"c�e��#�\�s����s��6n�n�wܼ�q�ͩ�|����;([m ���V2�8y�	��ɤ��ABZ��*�/�Q!بS\��7��K��B���l�)��
��u�N6��ތPVk�f����Jdc��c��2 �=�����K�.�@_c�ܕs�n̓Z�%}e�b�B�2Gae�ѹ��_fdv���ˌNOb-/�tɯ���|���u��78�n��c�MO1�8���v,L�ci����l�����UFg/1t�4C��1���:s���Y����Q.^��W�/N_���2�2u���'HOOS����iĊ�\���9m�hfK�X��E�d�a��h�iO���}���:u�c�r�[��5��$�VA$��|����\@U��@_��W�������~�����'s��9�(ƶm676�tډE�e�,�,s��)��ռ�]������[������C"UA�E`���!AH!q�ν|����x*h���AZ�IEMQ!�(�GY�@%t;r��9�����Cކr
Jc޿��{��x���o9z����9��Y��F�M|=d>0���i�RAH�����
)U�h*q�T�e
H���BO�@Gh�F$%h*FJA���R�ԦN�y
�U���s�5{)��8v�n~�-w��W���b�5Ûo均�����ワ=���i�8�DA$� ��&Q-Ab��UT2�P�@�|}�L��o���'�(��(K5���fj��:rjkz��a��x��vym�A�x����,k�g�/6���y%��dN��Wcɫеa�o⦡ElV�zɧ��YҮG^B.�)��\ǥ�(��urq�~|&Tɞ�c�����2�g(�O1�^c��d�w�b��.��.#A�P2C��RCR^���1���u髴驶�v(�:����6��&��.E�@R�+ce�8�@Ŷ�GH�AS\�9���5=J������y�E��s�_x�;�}p;�$��1�aH���u��]����0Y[_�7�w8u�Q#��������/�:��R�L�M�l�.%�뱼�����}~�C����������jR,TU_�e2 �H��ĊDc�!F�%	�碷]���GQ͢t4l2�d0d
|���a����R�xL>�8,���>��{8�s/7L��_|o��fԠM�hs�?G��'����Y}�8յe�l�^�L�"D��ؠb$�]��4"�n@�ӂ(N�� R�(��ek("��[�Y;�3�k��u����i؜��"�m�j�a���<�8����S�6.�����7081���ĩ�,��@ر�B�qL(��B�[I�46AF�����!gP�ۤ̈��Lme�(�P4C�f�T&��[S�dM��A�x�&�� ����=.u�\U�(]^
�LV=�b�Wa~Vay	�V`���M��^�Yh��U����}kH�(@�DfD���X[�PYc�������m��|�?K���Lt	F,p��A`K�T�cKM"��)�q�6K�j"	��	z�u���0�Dy'Á�	
�HE!:	�[7�uh?}� ������&��w����o~սܴ�(3��(�'�'�B�T��m������(l������'���?~UMj�ؽkǎ���������4�M�H*��177�����z���������������r��~D���!���_����1&1va!j��!Y(�X�kTs�u$(>�@Z�3Ub�����e<����Tu�j��v1Q���w�ʽ����fd��ӓ�bOҮ9q���+8Rg_� ~��%~)�T��A�#:�h�	B!���"�@���R��(
BU����������$XX��
d{�)p����9�/��\��Z���t[qؾc7o��m�~�,�#{��#����
�r������JD�k�SH9���"ȩ��*q؅v4�~_2\�P�ܚ�b�0�a�"dL�ԋ�ˑ�f1l���"[.�*�sT;�TMPWکn.O�ɣ�T�AZ6�v��J��g��=�)�H��fɬ�����f2	ad�b��v���A1
��WFk�����BQ�(Y�`a�RIf�da�4T"|<�AlK|bSŷ����Z\���)i��Q���3���.�]Y�<3Mq�M�YK�R>h��Q/�cV$H�����c��^qGn<L:�?Iya2�h�6##�4�-4U�9�;�cf�fy��@�P��i����P2�����ĉ�pl��{�����t�c�⟪P.��lV�bə3�X^Y�u�{=x�����Wb[6�h2�B�Bk*e���IEQ$�L��� N�貑d��h�L��2�W����;i�γ��#`��0��7o����	�h�~��=�,M�f��ҿk��v��b&������H�VE�U�m�Ċ�A"V%qc
�! ׅ�Ǵ�-��ϹvIY�8�e�~��b0l:2@S��#Z�B(���3��;8;�"���5Xf��6�m��Αavo�MԔ�q��9����1��BU6�5����05��u�]��ry����ۗd�29pCD�e�~�F��
�H!��Ė��*�mi*��BU4�a��4�i:DR'V&��. Si�T���#�%L�f��a�{ɏ�DJ�=�<�k8+���2A��B���tu��I�������MVhR� �Y��6u���L
ٗ��E�WE��E+�q
��i�A�/K�����@8X �K��YDu(�>Z�-��{S�R����k�6kXn@�Bȱ�S���eZ�6'�.��Fyūn�w�?��a��>�B:��R�ն���(
=�v�@7T���yKT]�_����'x�{�û~�W��_�%�0D��\Z�E>W ��p��9��.�_<���{1���|�x �1)�P�)����u��eHDa��[`���P�)h�������,��P�4Z�P[[�������B��.�>���t����a3,sҕ4�4��-<�⋼�7��=wS�>ae��٫TB���UH� F34PDB�"�)#�s�(bni=�:��J%�	�P�~�\Y�5;d�UjD�!��t��F�ԅ��#R�<{�
�8�];�[o��8��N��+�Ɏs��k��B�K3~�Xhu:�� �2�<���",��ًl�x���F�BL ���.��*�	J:CWQi�F��k�H:�O�t�[t�m�^ߐ(�����%�d*>v��`=�R�B"`�
VJ'�5��.���u��YR~� �y�@.�e���f��m�!��
ŖOΗ��_�W��6�\Y�䅅u�[�之-N�5�����J�3U^�kq|�É�/]]���O,uxr�œs-������-��m��t��g�<q��s�.�\��!���%���	4	�A�,����y]�Ȓ���{ٹ}���˘��%�k�!���*��7)�;���,,,�7�7��1����o?�9�&q�n')�l=j~��ޚI�4M��}�e���&/�>���<���ٵ�r�-(B%�BU��E�ؚT�5�o�("pb2���yZ?���y8y�����t���!e���8��}�{?Gn���v���s��eOI��~����?y��]��|�w�J�/�>�,/��-���D���#T�a�j`*
Q�BFx~;9� ��DD,Bb$�����A!lq>���:�S90ڐ	�7QjW+��-�t	�V���7S_�c���M�z��ܾg?c}�\lR����.��m�>;��U����`t������J�fq����\Ai{4{�Y��M�������u�2Ý���0S�n����xvd7O���O�Gyi� Ofv���>.�?Lu|�h�v���;t��툣wѾ�.�׼����X��8F��D<7��	!N��2V��f��*(�yF}�hv��TQ��H$ڍNJeMUXoEDy�d�r�,�d'���zM�F��h�4��ͧ�E�ZJG�?��p��g� �\�F��s4�6T��H�i����x.cp�d��&o����2����1��&��Ւ���Cd�)�����HU�I�����*Q�뉪����|�`xh�0ٷo�_��{E�׽�u>|-���k_�:����q�V�Da�e���I�$u�͍uf��(沘��w��n��F\?"@C5->"\B�!"G�A����Q��v���!�4j* �(�A5���q�6lC���)�ۿ|��̷�F%NϺ��#Cq{��w���E�(u�:}��kM��A[@h����c뤕/�`�:�(�$�:�l�� ?�VL��	������膎!>`1�%��F��� �nr��"S���.Ƌ�c����ef���(�cL��?|�>�mz�V�K�'�7-���R�	�<�@?d������5�f(t����,��|����F�7�xpv��nVx���|�K���A��Y'�|����=ln��lo/�fs�>V
%�c8���+xh��7�W9-��V�m�2³¼�LA�Q.��\m���J�@*2��V�%�u�:��51�wi�:A>�(g�x����C���G�)���#y�(W�=<H�����V�G;|��v
�����^O�{pŻ�0�ͷ���h|7���4R��7L������22����KF�ƇĴL�<Y�I��a�6�?����8y�$�s���?~���a�&PU��~T5��q����>��qs��M,,,p͡k���/y��o$����Ip!�	|7h4��+U*k��۷�����,�X_�L&C�U�� @EUtTb�E�T]Iz�~��r �C�S���`�A���.VZ݆��O���4f�dm�2ii�c|���_�G�=Ho�ē/���[����I�������̓�AJZ]?�7tUōc!�MCW��0��l'�u�V����#)�H��q�P�8�\�%�	d�]!E����\�?�"X��O�3���|�w���3��(R�<��	�Z��}7C89�H�B�}��S��T�$m��HY�Q z
����*2����Bm�sY���؄f���,�3:�n&M7�&Jg�Uh�*'ڛ�E�ˋ�B�J�e4Bţ�h3��l7P�F�/�1��7�u���`ծЕi�~��b�f���ca��k#Jzb�*�e2�x��v��'��,�� �4�z�A�<A�ج��KE4O�S4��	^��I���Ȥ�
�zR��:�v���6$U����*c�]��{�M��v<�A�v�c�����9YxMI��r��>
����';����)�q́�����_I�S躎��ضM�z�DQ���g��ٳ���!EQd`` �HmQ��*&�8&�N�hU!�L�w�7k���EŴ�mr�,�s-���&5dRS�L�F�B!��d�$R ��6���Pi�1�J��P�kAY�\q�:~����FXvh.����s���o~������s�տʵ�"�3u��.{�YU.�U]f����][��44M#��0"d	ÐHM�U1E� �D#�?�@"�BC�A♈cP���F���nH�Cd�nAc�c�m��©��a*aDe��\nq9;�N�����>��;�|�
��:D&�!7h e��nM�[��l��3�$�V�Ē��R~��j��y�v��&M�{��YXd|x�����J�r�����b������|�����=�PH[)��6�����Y�mR ,�gm��|�o���	���d�Ҡ3<@��~���(D��.����d�l��i��<����U��6a��m�(ՔC�11
):�D&��5=�J��>�?9�O`5T�L�{���n���jZ�:�㣬E1c��8��O�r�\�?��?%�ˢ��lb����"�e"D�U��[X�t���c;v�?�bdD1�碘:�lY��$���:IaKxE��� �����Vd/CVWW���h�����Tj�C �'^�
cc#4j5�Q#Օ%��az�<��N�X
��'6�Kۭ�
�%�T!FC!NeA���Ϗ�b�c���!��a��T��O��k�c(�|���+��~f����/������x�gp[m�.O�+�}�+�ɹ���l�v����D؆��*t�]T��kEH�@�a�� �A2q
E��nҍ9*�������t��0<-��˛LMN�{�~���k�x-,O��k'�7�Ǿ�!�Wg�//�E^��_�_�-C~�T�"B�䕀!�_��=j�*�c��q[��������n�n�q[<��(��mz�9
�M�ΰy�4yY�ۼ�P�f�/���%���鋧��x��B9rY����2��:�*Ks�36Z�u���j#c��}��3��<�u�\j��J�V�}�n�����b��Y�����g�|�	���w9��Ӽ|�&�����x����y����ԓ|���+_����������_B"�k�QQ�n����4�#��,�묶k�x��Da�Gn��G&�7AF�&�G0�g��c�l�-��s�K%�fmh��cR�C,�FWT�� hu�	n�������c���&����baaqK��}����k_����7�ԧ>�����w�/~�|��_������~��~��?_ܡ�>B�%,�feu�0Lv���Y^�����
�F6G5����S��q����%:2��P>A���!6q:���T�S0�C�+�,o������sԭ	��m<v=~볼��x���ObgC��.���ٗ.��܆T���A�q@w�Z"*a�4|��	� �4�ƴD�q���խ��gI>�1H��V�l���
v)�26�U�\J��^����Fѱ��{��������y�[^��7܊��+_w�����*�#oQ� ��GJ�}t����&o<ˁ�))���]|ׅ0$��0R�!�J17}��<��`������l+q�M�������o���ś��Z�z��x��s��}��1����{2,N���ö�~F�%��f���tZ!��XoET6��M(L����}�$W<���<���Y�W��T6�;-��`��4�g�ѷ/��:?y�����?d���s�Lav6�L㮯�!���ۤM������K�Oq�;���na׵�����/�����Gw�QpC��Kj��yKeE������	_�J�wӼ�:6����=t�	3XW5T�\t�ďBTUK$Ł�������|�'�v���|B������$�����o��o�g��x�	������}����=�x㍼�}��ܹs��K�h��$&���w��Z����"W�N�[*!�aa��Q����n���&č�S�=��p\��N��t��5��i�JB&�v��4��V��F������L=���L��r��7q��)�����W��K'^�ʤ��w���$�_\�ªK](1�s�6ghu<UEG��q�t�0��rQ,4�H��f���>A����y]��H���咖aM���eM�3p`n���2���C�Pq�5�
)֚-N\�����*���bx�����SO]�[�����t,�D2Jb�F��B&N� 9&!�
En[5t�7*x����eb�vv�Qʦ�5A�?���F���Ncf��gΟ��KL/α��ȹجT�Ln:��������߆��`��Ⱦ���x���r��J�j+@��<Z���m\%`Q�9�����x���1�����.S;y�~���qj���M\���]w)컎7~􃔏��SGn��{^�z�� �i(XYM�2�շ�Cc�˝�}ۯ;­������ߧ�����gV���+@;R S(�ɡ�z�㄃;��ƻ1?�^�x?����m�pw�˪K���M�0�� 4���"Nĵ�Gy����?���|�j�J&��g�}�����O����o�U�zr���!���DQ��8|��@��d�L�X���묮.��Vj͢�QE )��jU6��H�o{=G?�!n��ʱ���\��qfw�mײ�ґ�Ch�I�6�ޕ'"Na�e�tT�BF��6��:��8�k�}�y���;_�����7�k�0��Sϟ�u>�W_���;|���^mB�(c��ڪ����G	�U���U�0�B��d�D��)�R*B
�B�P����J��j��7�v���M��M.�G���
�zz�M-�6r���o/��o���s��z?W����Gf����#^<1�u�+�s�6V׻dEՑ��Bp�
��'~FArT��(���'*�KK���m�����J�\$P��������c� ����_�^��W�˃��	?~�I~��'x��O��OO���s<����:|��_��Y��вN�Kgzu�9�F;
��:H� J���@�V��B�g_|�����e�<6Ja�����J��++4m���*�.�VY$�ҹ��7������
_���yfy����^,P�$����$��c��%�+W.p��V�<��s�:��[_�
¢BS�A(PB�7?�r���Ɇ����^��o~7���s������7��wi&~�P���-U��v	�)��&��o_���}?�3�=w� 	��t:���lrL�^�a!H��|�S�b���|��_%�c2�Qm���� 1����Y��D54�^�����f�ȍ�փ?��_zՅe}�֊�կy�� l��F����q�"}����ӉQD���)�5��V	m�����ŗ�g���ι'���>����y�b���;�q���<t�K�R���k�dp�(���P�(R%�c�hB!"��'��V;�(LRya�7�I�BE!ix!�n�H7(:�m�t�XAL*�p\�+.ͪ���ğ���G��7�����"�:e�/�\Y����E��ФT�͑����]Y_�bլ�"�%�`�P�"�P�[�Q��U�}|-	����4�mV�*���33����&>=׏�Bճ��ԙ��J��v3���1�4v*�P^>w�.r��W��J��B�2ye���EV�W��h�!?`y}#���
q&���mU*��9T��gxy�jN�ԅ38v����3�{û�s��o��-w���Q�(�D���L���R��+_�j��{��*?�Z��%���_��65˙'���n������Q�~�=\�-��껙��H�H���!j��Ų<Z��n�Lc�ir�<7��Î����퀮��	�^���ΐʤ��6Y^Y��o�\�ȟ��'�ηD�*Qr�-��.?�0O=���y�G��˲�V�|�ӟ敯|%��#�@�윱L�ު�m�Rb�3���"#�c�H�6�V��f����g����Ɨ��?~���;<��i:~D�@�b5	]H4.� "@$HUE�|��.��Cδ8u�2cC�|׫��W��Qn����֏�%�>Q�K�5�{��ήpi��>���odp�v�]��?� =�5�̳�QRd�+�A
[�rE�I[1NT���*�FB!VZ6E�� ��vCz8�JЊ�C�+Oj��Vy՛���==�?_���CE�m̱�lս��\ǲT�4��*���kT����@����7��DJ��D�h:BUq��n�P�u���9Ο8M�Z�ؑ#���������� WgV��z"�L����	��$ĪJ��nڮ����ȟ��O��b/�8���W/MKp#/�hD�'D�a�HM%�N*�]���-۷����n���%���m�0/�~������9p�(�у��`�ĺ���_��י���ON�hK+d5� b�V�v��+�m%J>�� ���
�@e�(lce��5��Y�L�M�������W��M/�j�it����"�Q�H���i��?�"������=��1�W�b�&R�_��_�s�N�����_�z\�EUU��6����9v����x�������SPԤf�eN3�hk�ŶSd3|�G�Za�V�=��N�|��S�\�:˹�S�!�o�al|�B��;��@���K+�]Z��h�<W��)f�wB��.�����ѳ�闟�t������?y�
�}���Q���w���mc��p���e���Q��#TEA�tM#��0 
%8)�0 ݤS"A��$� pY�\e�Ra�o�&�[u�@)�@�¬�6"�4��8��y�G���￝��װ��;H��js^���#�����"5C%��2T1����v[�$�K:�b��
���*ii�Qz�=vK��,Vy��/MM��ui	H����d{��(l��N:f���ԖbΝZ��f.�u%#�~�V��1l-a�����j:�J[� ��
�b�E��c�QF��0�����Cf�뤳e����5��`�y˽7���o<%$C�6WXݜg�7K1-�U�x��(	�q���.��V�X]���iP��X��R��&{����E'n���t��d��a�/��A����e��3Ϟ!�x�J���(�DB�($��6	�����:�P�m�?�ԇ��C�.�\�n�epp�r����0~~Ǽ��{���?̅��׿��K��($�h6; 5n{�mAD��'��l;E�٢l94��X�:M���x��Ǖy��X����båA��j(54���*��[C���8�`#,b�#��=d�!O���dw/�7�'�������a�A8����o�_��^1�ՍS��<O�̓�Kf��0QcA$$�0�����*���E�H��Y	�O��V@�U�nķ�\^u)R�/ΒJHw0�m�x߉YT����+�
����2Qe�s�ϒ�7�瘮��Z]�76���std���Qڣ��n`GP5*�`���F[n���S�;�G��(!J��Ze�m�Ʋ(�NN�`��V_Mh�R���m�\�{?�\�\:̀�0�z���~��C ����FOi�}��eT��t[�7a��g��&�_���h��Be���~�[8᯳��G�����#?��g�g��"����g�zX��1={	]/P��1�d�4����V��r��0����y�ß��w��݌�Yڎ�;G:W�/W�?;DJ/�7�Tg�f�S�wqt��F&�AfsLW7y�����o��COr���/\bU��6*-���}����`�K������o�k��Ot�,�c�n����v;�ZM��������>��(bll��}η�����_�/��2���������)d����쓏�����اծ�͘��ۖ�-�U7���o�s��,�t�צ��Z"]!.�[Z?��j�_����i�+)RF�[Gu��o�T��VXX��w�M_�L�`��;&��o�t��2_c킏S�l��iR#T�[�ȲŊ��"R���܀��Ҩ���A�y���!	Q?�я}\pf~����Ďm̮U1�9�HԺK�Q��|��!J)ĺA���)DJ�p,��6܃�m��.��~�J"�b:����7Q�-*�.b������i�S�,0,@�1��NP�2{�!�E��B֛8ݘ@5Q"PuU�)�e��蘬�-c�)�T�Ø�F�V�E��MS�9izzJd�y4;��*X�M_/���Q�$�ae��^q��NR\����v��g����{�K���η݅�0E�� ��Jwi���Q+���J��F��fQ����y�Lh�{O���&�W��կg��Y>�r3�����Ϟ?������:tǤ�ma�
��A�ea�,k���Xq�u;ĵ.E-�唙ku�ǆY�hQ0N=�/�����/�.=�l+��N9D�������$E=ֹ��ױ{�n2�aQ.���_x;�|EQ��[y�+^�7������K���eY���p��FFF�,��B�	���y�|�I�0I�:mL;E6�f|�6�h���ҋ/��1;�A��J4CExk���Wp���0�>K{�dE/BT�t
#�D� 5F��hQ��~�#L:�$B�
6XJDNˡI�y������w�b��=��1��IWs!�(����	b+P)��4�{J)�'�B�E��s���kK��;�2�x;�����G?���aja�f"�a�[���YZ��DϗM���@��vh
���L����BZ2�:�`��Ie
=%:��"#���!T�"0E�)$���>�m(D�d���2~���I."�v
�-��Wf��t�xj�������Kk�/lP_�R_��6����
�n��hҨ4Y��$�x�.�0D�թ��������2��&�Z�V����,�Ks̮-���w��y��nc���(+�ȍ&J>Ϧ���U4.���?�-���6[����O]"�֙�ڰ0Go�M�Tؖ΢���Իl�x���%][g�rk��Z�t˝�&�r��'p�S�=�\^x�n�a����� �ҹp��v���^B���g�f��%ƭ<F�A���}�Z-�g���<}��������՘���-��d'c��ڨ���k	SY�0����a����1դ��:��`�F�Hߊ��,o��;���4�M�!���ؕ+�<��O�5۱P���z�>ι�g)��(HV���1`I�&Z�"��*X���O^@��:q+�"�@�B�(9�X�!n���)eHW��A䋄!������w*�NDʴ�-zT�1JJ!-}:fUF��GHK�󓑶�b`oHO��[4�.Ƌ�&�v�TW���x�]�^~�sg'9t�D���������J���NQ;
��pS����w�=���ֹc}�k��Z�ed�"����W��֨�?�����:�UV�*T�^�\���TY�\ǯ��Yۤժ��v�f<��ݸNh�X�2=�4y9MGmkDUrY�:�[�c$ޠ?��5��+�F�lv�L�kTE��p;m�5dA'h6�� �됱�(�Yk�סfJV���"+ºG��`jc�y%��j�$wdF0�g���7q�䓈�e2�4���X��u�V�i>r�r�E�T�4�S�p�MM	pۛQ�`�*)b���N�P�):a��N��9�Ҽ�������)��Na{H��g}�e��w�{8|�&��)�ƶj�
ٴ�3?�͙���Fge�t��b��Gq;T�L��[`dm�}��*v�m���{��,�r�t�AF!�T���xmEU�U��;���uR�4�m�����?N����|&''q]�b���y���?����Gᩧ��S�����cphMQX_���G'�r�L��s�ئCoOr=w��_����X��g�l[�'sy
��$��K�Wg�<yۗD� �}z
O� -Њy�P�̃�V��)hmV�;�jd�*)RV^���!XK���*Y�P�J�~�i+K=eRI��
Aղi	IS7"��˰d���"ܔƾ~(���^����{��t�Mr��G9����+���(BDk���'(b�5���� �Bm]6pe��IZ�\
i���&nA�&Ik>��i��:>�������0�A�x���D��D4]B�b��U�z/��u������r��y���2�{�>Y'�e;H���e���/e���UP�e��1��'V�(B3Z��N C,��"�4�֛EA�0S���W�VT�l�+EM���A��݈�	�k��}��}���L�����Thw7�#�7��G��������c�z�_��B�?K��L_)�*]7"vL���@�HxYZ���������>ζ\Bp��3�/������<~��opd�8�v��S�_�E~4y�v�N+PP��PC���N+�$�@��46���,����;��|�e%v!M,�24��w���|���u>�����O����\���1,ˢ���}�C�w�}�����*��z+���J����W���Zv�ڕTh�]�i6��j-<@.�G3t���+d�)�PR�T�t���E��Y��tT|?&,ݦ�A���*��h��	��A�(a�Y��)��3�]�v
��3�U1بm0�ۄ�Jl;��Y�2�Hc�FS2K�~U倗�2:��gȲ~�����6����EǢD����
�>Dxˍ��2�:B��ں�Ғ��I�Zpx�j��.p��Y�ZA2R���XxR M�����FD"��b��"�zKU�D`D!m���@	����X��>�L���e�k�eڡJ%Z����΢�ơ�܋S4^8���oAn��-�p��&����bi*���������R�n�h��P,����SxRŴ-Mcbd�;���B���_��ow�pZm�D�0���3~�Z��ǄG��@�v1L�F�b�-��]��7~L�R`V�\�oaiw�<��Ъ0�1h�K��b.>����"M;�;��������]-b�~�7~�� �h�;\9���曟�=s��|�3��w�7Ӡ�±�ĕ4<rw�ǃ]���s�m��{>��Q�E%����G��8�}}��}������(��忼�(� *@տJ����,��ԧ��'?��Ԑ��(�x��y��^ǹs�ػw/A`�:'��̇���t�>���j{����11����dR�==<���l�x��{�Ԗ��Q��]\E��٬�	=����8̹��<�yP�Cw����on�L4��� �E���@h=
����لBC���'-�� P�aj������>�*�t����S�|�!ٜå�e��n�ݰ:�`KҠ���ދ�i!���9���?t����d7��xUdB*5�EE�`���s�D�GD#l U�f  ����Q���ej��ED�q���Z�f&��X8�q��Ȇ��A���u1�keh���w`��M����aq�7n�F���N�奫���z��_!����z�ٳQdD��`�;&"0U�N����s��;��)��<��|���<�߰�O���	f���	��(mUp�_}#���2��/c���a��V�9��gS/N�BE�Ɇ
��� �#��/�ub�N�_��~�|�ce�>�~���g>͟�ۿ`(.��1֟'�m�����L�ɣh��:r=��D}�B~76u�L60���ZDM�AD4}h� R�(�ŅJH0�F��)m�b�z���	}=y��MN�t�w��F�"p�;ﾛ�����^�zRiM�x�'��׾Ɵ��R*��p$	��?��Ї�z�*cccDQ���c��(L�Լ���@?B�F�JE��w���(hB��	�B55M8���A���t�1��KQ�F?�T�)V9� y���Id���	`+p����](�Y_'���J�3+�JYo#Z�&G���D�.
=q	i"L(:`W�tIh�I�F��K!Kp᫼��bɤ������+h�$�l֦iU]���T"�a�J ���[Y2���Ү���.P?3K������f��=���C��a��&�cl�f2:M�.O���C��<�0�Ne�MV��^ڣ+��-'E��m4/�%�n"WB;˒�g�^ºO.t���3�}�{��Jn>v��O=�ȎC<��z�b�����i<5��P.�u���D�B-��Θ��կ'
%�����]��K���.�����|�_�si�F&�!��x��]����	�����j�����[�\��`)C��$�������[?�9ס���^��W>¹/�d�4CGob�o~�ϟ좎�'�Ǐ~���k��p��ny�7��Б>��6���_�7�m�_#�&� ��
(͈�f�J�na	Ev��\����v�`uu��e��\�Hl#�s�"G\�z�'�5�n�K�@�F�Q������I~�����R�D�?��<y�$o~�r�
۶m#�>���(�$�IQ(���U�B!K�Zg�V��/�l4��tg�8YU`W|L_�**
j/���(���i%]�(�VH�=A�s�'Gl���q�U��"fc�'j�0����������Emq����	�����d21�'NR�a�}�sq�$�o������9��u6�^!_�ax�v�j�3��W��
娉�&�[��M�������I�F���P?��\��N�������Rh�'�#2�8n����և(::��N�����W�^_b���ldT��/�G&7��-t�q����v����B��Cô�*02�`��̥5�F�`�����0���\�M���Q�N��{���Rv��#\�e���;o�J�d>7�d�#�}���>�]|�eF����s�(�е�Z�񆮣ѿ�z�*��T��>r���=x��J�7񵗗��爷f�gs�	��^�^����k���������^��xf>�Wu�a���8����&�obz�-\>̙���]{7�{��c���G8۳�;9�Q���Gtݵ��j�����=���?>�F��q&H�1������;ވ�Ʌ��w�Q^�;fs�YǶ���c<��_"t�Xi�n�I\M����wږCi�!ֽ���B�ؙ4^��ł0��Qm��ǝw����0M��x���y�[�J,%�}����/�cc�X__��'�dhh�0���k_�Z^��W����Ų,d�n���7�E�Ѣ\�ann���~��G�\.bfs�w�5j��M)����@�j��,�f$��!b4�yu��&Nm�be�|}��_�� x!��\����V���_�����������6z�{��:K�v����d��Gi7dE�}��ǃhk�����.p��אS���N2ˡJHE�8[�-In�E��� ���SA�bvh���G���P���t4�&�Ѷ���_���q�D��[�woG���I�T�c��*�,<��P�)���/aDu&O���z��0�;BE)ru�9���h
%=bZ �iѓ2��\������i�j:�!�8|n�������&n7`%��Y�Y���_�˝�%�L�G7`�+�Өm�uR4;lӡ�{ĺ�/-����=H��d8�*���9��%�� ,�׿��>�{~	֫|�[3p�]��'�A�:�x ���4ddY����Y�C>��Y��P"@�y��axj-����.��+�JJ�-���0x<V4>]]�n��t�������ocq�n�!0mS<��Z�BG��m!�D�:~����*����(P0t=��Qerz;�fee}��rij��{�`l�ST]%�ɢ(��������97�x#�mS.����@�u�������{�瞄{���q�m8��x�mcqq���Q���	��B�H[*�(&\���*����)�
�!	�B(c���#D�ƒ\a!��4U�|���=Ɏ3���`]������A�7����]N`�v�а�WUV_8��-�.��\8��)ts=�ݶ�L_?g��S���u�`��)��%Դķ z�aIU@��2jѫ0|(9�T�6Z.E�:�>	��M��
}����g�B%R�z
C蔍,}v�8�
dK1����Q��m�s��q̌�d����2��,W����ڟ�ކ�"�C=5J�(�l�\czTҰ�6��]�K�>�K�o�n/S�}HK&�.K����b6ϔm�a��FK�Y� #Ҫ�f�M�D	��� ��|]r#�|7���m��×�t@)���b�A�ȺС�2�.P�02562P�o����A�_�<Q�4��l��I����@=�ݳ6Hr���\���ڤ��iv�tb[���(�sN�>��u��j�hY쮎--2����&��ra�
+k��.PY^e~n�=���W��o���<�Џ����o��o$�_��w��W��j��ů�+����ٟ��b�8�y�k^C�|����s����;�C*�"�c��#��|M��(��m[�=}��ېBA��@CS@Sb4���s�L�N���+�8��"�(D#FCA����w:Se��&^m	��Ѣ�j2��6�
A9�"�!��X�����X�����bѳ�0�^{?���V�H��-���Cۄ5]�Q�kkB�-��� PTd �P�5٥w�U�X.Z �0F�e��;Y0��^�d\�)���+E�f�L��� F4�f�W(w�i,���b�;����x�ʩ6��-t3��&��-��
V�_G���yI.ǐ����C*���8&t:�J]�T��LG���R��cI)�����t�$,Rx� �iЫ��*����KA�Bc���w]�eB-�VA�x�Rm��a$;mPŒr�GFUɵ}T2u�r���gGܡ�+)F5"+�)=z�V-&#GQA�}�n���[��~�������B;f-(pn�˝��6ח��:Q�ȭcZ-���W%�
�Hv]$k�)Ad�L���v}z�,��
�+�L7�9[�䱳�t׹��#����/�_�K��E���Wٵs7qc[6o��>��+�B6��G��;３0���a����w�����)���>����G	�2�FX��`� ��s�ݵ���O��e1�r��bk�Xb��H�"IN�L�ժ�iW@���~6���@O
�t���Q i�g��pJ�h�C����� �KO���@�X�P�۔�Y���PT"�EI{��1Й�p��?�?8��O�����7s�2�R#l� � �(ɣ��>��@��G?�qS�{�<��a
�Pv����(��V٠��(�v_CE�1t�6v����~���%���nV�&n8�Ǭ<�}ܥ��c�2���C��m��m�]nP)�ba/'G��pD!,"����U�錆vH�*)C�33���)�v�L)O7h'���t#B��n��)��MWr1hqHKD�,����*
�A<��Q!_��jtY�8���K�FG�t;��jR�6"m��(��o�("�`�L�GD�豚�b�FD+���Y^�~���S�*U;E�P��yI"ǖX�@��
]B��D��5���-�"��|ㅧ���nN����� ��	�@�n,!V@*�X�Yu#�5�϶C8q�"�TQ��j�FGфB�L�Y�D15�;|�^qo�������j��!e�����e�Νd�YTU�y�6�@j����'#TB�'�#:n���S�2/\b����9s�V����	�?$�BF�6��
�0�'��Jt���粬n�C�Ĩ��Z'B_EUX��.��o��%38���ס���͔�6��� v��5w݂���0����=��Cv��ʱ��c�o�΍oJ�š7݋{�4��N����1��P@KT!�.YW��|���G?�:Sg��😱��Dݐ�^Diu�Z077I<8�=>N;�0�����e��ZM�}`���\z�I�+(�9b��֬�]9O�4Dǲj6���v	R06���䄊�vu�B�5X���2Y9q�ŋثU��u¬A����R詵�Iw�N%��T�'��[F,a��>��O�-BA!B!
W�y������&���æ�ؚ����@&�z1�0�\�8���~�?�u�8B�R��-o}���3����~D\k!u��@��WA�]�$~(p��фN͒}&�z��\������	��9qj]O� tE�@�R!�!�U:�J�ؔw��dr�{i�\_	7k�8��Ս�"�\��v�J�I���rl�WWPTA�ۡ��a��TU'��-N���>À��&�>M��]~��L/.���^���xy������UT�@M�W�3�l�q;� @�$���cU��f�lT0e�h����}.�XA�8ƑӅ��E6i��T6f9����_^'^[fu�*��oTY��gH�,��^С��Lj�F]����{�~�1��)�z�@�Э�N�Ħ $1��M3��]o&��7u��K���	a��0�I7��}��JDt�1:�>�5�������"�:I��q�+���XdX�Q�j�
��;��� �K(ϼ�9{g���!�/1LEjD�@S�d"��#��TU�fۅ�V`�'E'�	{���E�H�(2A����%���uE�I��PQC�@!D�1]�U����>�\�v�F����ɐ	u<[%pz�%���DU4���U�(���Z� HB&�QMӉeL�U�i��b�7:��
R!�)����A��*#7C5Fh:�b���t-�8��s�"���O����fO��9��ch��Adj�(�B�D8&���s�����7!N���2��B_*���2��Q�`����>����&�ٮ��v��(��x��*�l��(AB�R�h4�t��;]<�G
I�\8�g_x���aN�:���)�?t/
�U�Օ5lC����:����"N𒁒i1-҅��� o$�����X��\������T �����M/�?�8{����Fkv�e��5�\y�7�+GU�r�l˖dccc6p�&tC���n����@�&gl〱-˖e9)�*U��v�o^y�y~�������k����y�����c�<��r:+�į�E�]����v4�.P�!��uY�J2���x	��*�v�������=m��X��Yx�;0K�Q����?�jCv�5�?NS5�H�#+C���_��"�oQMA#�2� �iE.E�0���Q�'�l����l�M�����=o�%k�ak�N^��e�!\a���E%s6��Fk�$I`�G���3��ݴ:�����H�Q�-�OXXJaI��CU�u�U9�#�FV��ގ��Q6���+H�!X&[x��W�|�8�(����P����Uh�@Q��ڔ�EF���(��j�����R����O�X\D����>�0a[�5S�dQPY�\j���{�o?1C~�9�n���=��L2�n�f��Lw&�n��n����`j�I��`a��ٌ{;��1Gn9A�66V�B����p�.r�4#�$�ߧ�r��4g�2��FH)ɳ�4K���xL�e��}�2��'��._���㵗^e���s/!K���4��	�<Nq�E�W]iơQL0�nP]�%�
*�#��g}g��*1�~l�#D5/�ng��� À E�®
R��VcJpm	e��
�$ZU8�7yh�m��4�'�i+��4*T�ʠ�Z=[Z�-PN��oX���Q���?�C|�z�}�P�T�&R(A0�B�cMB��F����q7A�`�4RC��za�@3)m�㊲H	�9F�m�,?���n��7���EYA��T���:��;�Vؽg��xU>�ûYZ^�7�)ےx�D	���/�:fK�+����fu_��)�!��x��k���mی<�vY�G}�x9v���p=�D#���K�H\��z�+R
�uQ��	����t��f��d���R6�bq����E��'Z�g��A�F=m�vlZ����Cy4,���#�"�&�\Ń�W9܊�οB��9�$Fz�t�=���8�ǈ��#�,����9i��molq��AN�]cX�8�O��q���+XR���5;��vzTy�e�(˲H���(���a���n�4���"g4r��UΞ>����v�*�~�^��sa��}����VǶ�B�g�^֯��T�]Iƾ~�?@���,���"��am{��,k�4(s��|C@e��+nm:�`�zaj=#&Ca�\�B#��P�X[�g�s�5���?0���BR��W��HPu�
�#)Dm<۴B�y/fa��m��2�<�7\��_$H�b]�gn4eS����1���HDʵ)2p�:������B�	��q��;-�p�*�І���q;�0�n���v4�b��U����}Re5�hn�i� 9�ONqy�I�n��;HP�Ɩ�BZ�҆R�V�����<�i��q�,v`�!�����U>���(p�Yllm���FD��B�� �TTTyI4I�K**yU ,�d�4>E<�3)RYx��V0N�)U�7����Fv���Z�S�M�Ӱ�(�HDc<���FW1w��_r�����q�2Q�B��Rbԍ�S#07���kSd)��8��|te���G�1�����p�ͬ�!�+���X�����v-�n7Q���,��6Ҷ�N#DHQ�T��C�0F�����zloos��i�_[#�S����LR�%���ezz���.�ԔUg�m�7������ֵ��hod�,�z_{�hm��B�m46iJ�������^�"Pt�x�A ��Z��,|e]W�����~�A'���K�MM'�6��%��d���4���Xa�Yk�{��G�n���x������ed��+o�Tx8��prR�~I߃��B�GH����u$S�tr*��A;�b|�
�%�����.��>^�G�S�s��"�\�q�� #���q�`Ғ<ɰ��V�q�R�I����Ɗ\�$F�,ͱ��p�V9�6E�
�� �[$���B�$YJ��Ҍ�h�"��B˕\�t#E�'	Y�bʒ��%�c�$#�pC���h����~ׂbS�C�t��5C1J)�KW����f���5�Q�ب��<)�6�,&-0iN"�:�!4���X�׹��y+'�W�c�6�+(Z.Uӣ�\� @Mt�E3 L䒵L'"�r�al�j�KR�s��\�t�QY �n<$�LbT��ի\�v���k��l�q����N<�I��$������������˼���|����8��˻q����9T��r]�Ч�J�*cb~1Xey��򨋕�껩U�k#EŁ;����sX��2������q]���g��]K��0��)�?�HC.FJe�U��ـk��@`Q���FRHCn՟���X\�̭��6V}��[��z�����LTQ���K�+a��"]�������鴨m˖N�@a�o���r �@d!�Ω(�t#�<"C���6���wq�m?��b�}UG(*�P���Kz\�l��D�O�8(����)��Fi�(@�#Dlp�ǖ1L7}6/_�\��ؒM	����<�Ju�ȷ�q��i$N�ql%J
�g�W��M�(IȊ%,#ɓ��P��=��^��|z�bjan�`g�E�sh�"�ɪ�8�p\�P�4�MrLZ
<ai��ڀ��=��0�*C��%� !�lJ�p�!x��'��;}��k��)�,�Io�ۺ�A���P͐��)�N^`<��w{_�yS�qI��xǏ�,���S����r(�a@���hĠ�cbr�(��������(c�tͧJG	E��$1��E�����;r�ha��јF�ĵl��v�`}k)sS��=6�]f́�:��C�l�e,a���f(-����_�2v^�lA%ZH�e!�z�J��� NR�*�Siڮ�)�z�����J%��666��HZԐ4�(*[#��$�%%�c�����2�d�������_�s�}�|�g�V��W��$�����ꊏUW��UwmM�a�&��q�����ʂ���0`��Ud�F�F9ER(�L���lً�w�1�7`$!*mR6��Z�&�lD�e���^�T�C\B7˱,�JQJb{>���Xl�~�������N���"V���$���B[�б	&�����Yi	h�^��B��K"�@�����K��q��~��'>Fo�*���eZ�$q�z�i��������E�y�[U�Fd^bI��Ylc�rd����PQ14��BW��l���:��ytO�L|�2=��!�&u|F2��m��$��A�Ȣ	Ls��j0T.]ۢgی�Gz0�X�ў�Ğ�8�&P.-?d�٠��J8�0�a��볱��x�Go�O��g���e#U��������L`{Q���z}B��EhI�q�2����n�kW�9w�-�����줬'9����٘ӗ�#*ȵ!����HZm�����YZ�߿f�[���Us�ҋ��)]�u��
���_�)$�1�$�T��m����:B�Ѹ�U ����Bjl�
RO�(`�m3��o��=�no�4*�>�V?�+43��U�Cg	e	N.i����[��k֬U�@/��ϲ ��� �$#[��0ׅ��$G�[���s����������l��-�iP���"5�݌��=Tq�']Μ9M/c�$��s���L��G�� �"��)N�n�]�~�)ү��_i6gZ|�A�Y��kS�С_�F�>�v���-�뾝0�����YT�A%H,S�hˣr-.���'~�1L���[މݙ�r#r�!���j�p�7$*���=E���ة�>�����2�K�����.�`'���S)'��km�=g��O�����#$��"�]3,;B�a�Qd��R���[���q�o���!�'h�)��Ρvb�DĎg���9~���c��LU�Q�����rl��"��p�H���2��U�m�yZW��>���V���B�x��t����p����"[�:����N���/��^@��2d)�e�U��I<��H
�=i�h��$iԤ|d{�ť���_g��e<���}v�K�-��s��{V��Th**Q#[�e�t�[J\%JT	��4u��,�Wj|�&���5�2	�986���1�2}�[�71ox��m9l?�1���K��T����������)��������<�\�ȫݺ^����IT��!D�h�xT��K���C�|�O����Ǌ�����l�TM"'d�6Szĕ�?��3����`g����d��q��� ;�$�㣶^gF��B����'8���=�uP!�r�7#vO��m��6NhH�I�t��W����3p��6�Y-���9��s���]��A�{_=}�)3����n��ݟ	�D��|��N�x2�+t�%���ڙ3�=���^������7�ڿ�ڼ�;��(��<L��=�Z�3�Fɒ�OdMR8����+_�GC�_���;����#sn{��kk���q�����9��p��._Xaj��`��D�ű�.��*��>���Ȅ`s�P ����&O�M�IbL�
�h�Nt�ŵ�]Y
ae�!���-B%��f0FW�a����x��9�'��^��o��<�R&�	]p�ɯ�4�`�6%�sm���F�e��뷟(3��"���E��RFZ�����q��0�\^����4�6j���%�4�y�m'x�����Ϙ}�(Z:BbɊR�����Eap0�7޳���DJ��JQ�9U�	��  ��D�����
^k,r��0��7��������Ν�x��`2�ɰL�HaX�ju�F��2T68��
�@���<р-1n��T�u�C
*Ua96���fɫ��Q䉷��	�t��E��J���ao��O�k��×_��!D6LD�(,,�f�xc���/�;s1�i`W	�l�z��ƕBB2�(�ﱙiL��B����ŧ>G������za���χЩ���mF�7XIzҘ��CbQ{x�$��N�k0:�>~���מ�
Cν�*W������L(ٻk�_�������#��d���	�>�3Wذ�,/�U1��4�d�I���Y�}��_dx�%�g^�q�-d�	�<�*���T�AK����;�i��dq�v��.�8ebj��$Ƅ!EAa���bP��#��1�YB�Xx�B	��;4''ɀ�QLb$�dH^fP�
�b�p0bn����؞�5!�!�{]6�,e�=hۢ[挍&�GLG��a�qؖ`��0��T���e����B�w[6m��s�����a۴''��!�n�no�5cڍ&:�y��S<x�>.}�i�K��D��%Gi�A*��)A�:��k%��w
)�����V�2�CQ`�JhMiæ�X|�}���RH,�pJ�[*\� ��v<
2עH!���Cр��*c aS���*��f�� AQѬ
�+�D�b��a2B{���l�4�p�x����y�b��o|�|����ܵ�壷��{�`��s�`�^X���K�?�)F/��)z��v� �0T 2������[%7VYy�1��'�덷�x�L�S��'�2�/D{	n���0Մ_`��O�y�%��m��*mdf��z6�c1kI�����`eu�է>'_�=�������0����\����7˝0� s�0-�ٯr��,//��Cˢ9Ѡ7A��on�h͞��pm��h�Is�2G'�8A��Q<�q�k��:�*�r\�!���ݝD������h{>�m119��j��X����:j16�D&hL4�Z�%�����Ěj���.͑�!��#n�și�RRX��@y>^���4ZZD�ɕ2���%[��LM!'��}����P�}�Y�4�W19�^�G���C`��IG#LY��)�V�F�1�o2�G��#�b��
�V�@���:ѢD��TP���0hB�c3�I;-+$�|�(�vp,�q7���)4��$(� *-k��������M��k$O~ǳ(�eeЕ�԰ �`5�OFwTC����8p'��a6�v��k��zr��m�)�\J�*�wJ��Qӷ'Y�>��y�k3Y���6��4���sTO~���-�����}��Y�����	fL�;ᰚ�@)��]#������%�	��]���-�m0�� M�u���ė.�|����p��spy/�D�#�m�>8���>?�-'���V�/G\�t��@��UiA��9�341��$g�S*���у4\��Z$*�쓟�3'	�/S�́���w����ŧ���>�̮	���;��9\������('�ޥ����h2�()�B�m���`�����Ӹ����X.�,A�%�l�0p��LM���d��F��̘��e����#�h�(鰴�H'lО��	B�F�əiJi1**�EEsv���{h�̠���)&���/��L�u�D�&SS\��B���|��C�h7'�����f�3�xQ�h�C�+ZS�g^{��6�c;bS R��vc)�4��]l!hNL1�\7���Q|�3�b�������Ҝ�w��k���;����q�\D���������s��3f�)��By�=︕���{h�|�~ӧ*G�q��%*��WiC�q6	�6Z0ׇ������K{Q?������%�S��|m�T�UTxZ`J�c M�o�h�m��>���;07ݎ�w��1�7݊5��h�M��Sg爛"
������\8��sl�ep�A��s�U�=}��ų���"�%z�4Xc>�����\���l�~��ܲ��#��-{I)�a@���vh�'Y^������k��É��{?T�n������g�g��[x��9��&��-2��di���ͷ�c��w�[	g�<K��<�s�vbv��	
WS����9�<���SJ7��k�S=������� *y߱Y~�w���WGC܉6��w=� O��p+�
����0�|aIv��4��l�#6/r@��V. _� ���fs�Mo�R����R�z�I�^��-�o���H�v���`u}�si�ZXB2��C���^�P�
׶���xD������YP�7K���:��-��;��1����~�YG�\���@f�v�����.���p�����������$�c��*�I�$�2��v��]V(e6[l��1B��]�f��_�S�Ŀ�)���˘�'+
B��O$���{8���O_ķ@(�m!٘t��:F��#4��F��S�t�xi/���4�݄�����(�=�1w�t��a�_,]Q�u�T�z8AZ��4Xx�;1���R�X���U=�d��]�y��I�����Wx����oe|��c�`����7�}���ވ}�~&�f��=�ozّ�N�'���, ]��Q�����)��`=M��u�x��0�ֽ3\x�t��/}��,ő����}�w���l����;����x�Fr�*6�F�!H	D��e!C��c��e(F|�ɧ������#qpw��9Ao�E~�W�Qr��|�s|鋟���&��u�����]��UIu�":+P8Y���\ �R�lQ�%ٙ��)�ӁF��(���G�����C�^[ßY�=w��ؕ��~�_��;�Y\��L�]%gǦщ�x�2`���}L��E�1�,�6�g3�<�������W��h3�n��m�����p<`0aD��ƤyI��\:{�˯�!t�i(�<!++�%I�:�X��wnoq��I��z��kװ�
_Y8E��十e���]	"�G^|��ϼ����������U������P��,$)�W�^[c��M�fآ���#��@�%UU��:������_>ď�؏�07G��Y��5]�I�L3Jr
]!HJ�R���.�7}G��O�>�K5�Ԃ�������WR{��u�����~��v���/p��e��eũ0Di�5��BP؀,A� i#��2f��S�WA�C'3�(w��]?�ʷ���}o眘��5��&�e3T1���l�e����6������}���2~���]��Nb����~���1#����6��4D-������Q��Y�^㑽n=��m)����o?�I67^���;|�w��w޷���<���vB��@��、X�َנ�3+:������7?��G4��y�;�)'�|Ǐ?@��aj����}�p�U^y}����N��a{�j�G;h�Q=�),�>��+7���������c��{g�7x��K���0����-n>���g���q��,A��o��sƣ����4�CӤ�����$�2*]�i5I��V����v����L�tx�Co$�|l�"�p���
G*������`*P��:�T4<�*!�ǵ0U=kS)��EUW/xڠ˜��#��P�o��q�x<�.a<��c����xEBC	�[���B����� ���X�[�$�P���òm����jw@��U�� t��r�u�"����vlT)�,�J��C�@�w7���ݬ��(��o���
����d1ɕW�_���v�;~g7��?a��4����^���)�ۿ��c��~g�Ϊ�I$�4�֍�hQ �D*�l��(�Q!���������Wv�?��k4�G�xx�EV�?�q�'g��O���~�S���ȓ���5��빍wם���`sv/��4N?�Nr,x�U�"������?�N���?��C��)FVD���9}�ǖw�����,�����垻&���<�}oy�#�N4Ƃ�����M�U*M�u�#�83��6�mWT;�|��g���'9n������|ȓ_���/�{���qs;,���	JWܘ�*A*���,v�í����"�&������_�{��s�������l`�<c3�{�Q��W�x���:̷���0�s��#�2�PR��rUUb|/��l���i��|�{��>�y���Bh<KQ�ӝI|�&�r|��!�h�P�~��K*�֨ʠ,�E���w�A��v����
'�Q�+��f1�l��`��@`S��\U�J
G���L�X��k<��.�C^��@�Ƒ�&�$����f��:��mR�)��m
]P�9JA3�h7|l%�l���E�t�q>���4"�ҧ�4�f�I]c;�MnCo���;�1��o_�ΙW�x���y��7q����-�S<���a����r�o{�]����禙g���g����I�S?ʋ{C����"�D:5P�J����惕���W�^|��vq*�V^�ٱi��'�w>��4F���>ؗ�����%�=�y֯����AKZ�.����l�~�&5e<-RT�ڨ˾]�)3M�>���Xk"���|3�	�� 
��Y�{��D��"�x����mN�t���v϶	�?��kD����7M����[I��?Ζ��q��=��.!�&�SL�["s�ހdeH�"�|ް���?�L�5������s���Y޿��W���{o��w���Ȕ�}�y(|��i��)��c���k��]h3F�#��.Ck��7�'o:ʣ�A�p�;ￏ��u��v4w�z�8�ן~Mq�ͷ��G��%._}ug�0�t���4�������V��/���,q���^a+�a�(J��8��}{�q�w�X.��>���خ�m�y�NFC� ��Z�ӓ�)�-�-IZ�YF<�j�	<m�H�晜���0Oa��x.�cs���0�(K���t�۸aD�њh4�x�â��M<S録�4�-�,E�UQ5#�e��.qUb�[��
G)�$a��Q�9��|緿��g�p��]<�̋t	UV�9³�Eɷ<x'g���A��o�V��.�b\������5�ͫl�y����}|iӽz�K�|��a�]w��8I4��SW��Ľ���}֞~��)�8�xlZ>Kozb�Ad%LBE�E���W<�^�;��n�����t��g���?�C��v�%q��w0qp�<x���5=g�p��'��<�*eׁ����L�s?վ���,�&�<�2��	�����.����ǐ~�{��f��~��_����sg�����x����-������|	  :�IDAT�Q^��U�m�@�.XE��B����m�T��.cN��{�o�����������|��(����f��5�������[�ç{��(�PR1LF䮩�	�"�3�`+j�i�*��s��-�8w�<��#���O>����_�{�5���;9t���Ϟ�g�x��=�"��z���n?v ʊC��a9q��y�8a���ZS`(�hv�y��)._���3gx�������������gģ'����˯s��N�9���g�ڐ�1a�IZj�iJeIv�l��RA�b0
�� ��������s��1�%�h��v\tZ!��ߛB�po4�6e�����/2�0�K�v�,��DZ�<OP�O9�ƤՌhD�0 K2��@[Z�H�"�%�+�eN<p��Uzۛ$�!������c��aB)$qw���[�\��kF��B����G%<q3�Q5���vs噏c�,6[�Y<���1�\�h́��F��������/�G�}��wA�s2uY���:���͒]�̈́�n�9�����j\��]�����.��n���1^?cY
^��_��'��F(�Λ�n�z�%SH�1�.p�ڐ2Xڽ���9�^:�p����dr�LH��[�>�91NY���p=D�����t��Ox�UK�p�X�^{����?������7���[���Q�q��z���#lw3��8|?#��I:�7��	�+5����kC�Y\��'���}�k������)N������=?������{�~��Mɥ�k��x���Pd�xM���-!T%0&�)C"�9h�Pns����|���~�����y�).�v9|\p���@23�#�˗�x��sYOJʢ���B���Ɛ��4��*���E�0�F+��ip��%�SK$IN���o��� ?���uT=C�MZ��k6�';�$%ä��l��N��ha[$iIe���ӔI�k���h;6xq��|��p=a�T��rh9-�!O�5"��иTah+�P"$�Θ��hK|�i��(�"CP�	�e1=զ�h��UQ�{!P�7�P��fk��'��;�� ���8|��K�	'�ui����_�����s���]{ز��E�Q&�7��V|��}9bmS|�8��ͮـ����1SX,��d0!6 � ��I����)Va�&;���̾�:Ǹ�~��Y�?�1ė�6�=�Nk�QsA��
�;6���N�ѷ-zB-t8����	�Ԝo����fD8{��$��4dB�(&}X����O��}��}��u���u7/O�P�bsm�����O���z��f��~�<��yp:�h��v���i�L��r��s�Z1�%��������8�j�O<�5�X�ⵕ�LM�|��i6,޺�9�����s���SDM�AA� ]䠠�nb��v�Y�k��<�ξ��������{��M�	�ݟ|���?~�/���~�m��{����!�h��~����6i�יo-s~T���fmʼ�*!mZ��B�6JJ	RB�IV�m�W'1�m8.��x-<;$/�2����?��H�m��
�$#�"l壄"M���%�*1��q<BW��­�%��
�,�LǤnN"
��RXc���� �<l��FKK2(�T�@��)�y�v��ag��	j�#����0��k9�~}�"R�(�e0�q�!,��pQ���h��qa�c���]���ۜ�����o��4�ߌ'n���A;"�4UL�PZ8ck�n�=�+�A����޻r`����Gފs�v�&����R���`8(2�b��;���� ��
g��%v5��mw!�3�*����,0Ja��r�lI)�@ڸ�b�uظzˆ��ɤ`��]�D�����l�������&o}����Af����[js�}GQ~�SϽƾ�7��+�q}+���_aSN�f���"��Eu�X�`h�a��LC2��!�^��~�_3��L���w��7�u'�:b����<��
s��m�zu�R�_�kMS��u1��ӷ��k��c�����6?�ѯ�/�ȁA�oy���7������]�\<{�������^�k/��_?�X�h9F���=�,cW�!
2��9yQ�3R%�6#�<�F���:��0B`��롐�/,Ј��g�^����Ҷ	|�\�D�E��0��ʢ�V
����4������cҪD]T�BKY�@��ǲі��-*mR!�Ĳ���DH�P�d������ /Z,���|��5��R��#&�&����ݙ@��ԗ�yU09�"�|&�&8t� �V�
A��x�ǁ7=ī'/q�����z�@�,�=�;9��������L/.4[ע*%���I�����s��ϱ�R�ES��>�h��2�i�B�uƭq[h-j�`9�� ��x3��]�vH�q�0�k݂�����ia�IAbK�@�D��\4
B�0�C����Ao]��(\�������?�%g��2i�ʰ���헾o��p�0�?u��WzL����	��VWQ�˜���#�#ߵȳ�.��$s�w�5�b�6�@:
*CQh��fs�<��b(<~�c������~/k��h`�����{?��pמI�i�sg���3��=G���#N
66SD僊�k�pɰ(q��9Ͱ	K�A{�����O��Z���WH%�V�M�m~��������ғ_�{�������3%�,�w�.���o��y�����녨+()�\�ű=�õ"ۡ,*,)�V�0���`vf���%v��Mtc�I�(%NFY��+l�C)�
�m�n`=�#�3Fc�F���řL!���#7B�.B+��q�Dص�ڒ
e�����B`L�W+���H�t�FT`a�X��<�zp�����0
�����O�slƃ!R	\eљ�Xׁxs���w�G�A���c��z��Ӟ��u}��F!A�M��C�
���2T�Dd^���a�\x��(2�^�z4��� �U�9lU#V�H�M%$BhȮQi��%�I�ӯ<G�z���s����n'lblW��X*Ķ����!naN�@�m�St�7�Pd���!�D�3)1��1���6Ѕ]f�/|c�?~����0?���|��6�����|���6h�W�0�m�C�����	�T�3��u���V��1y���h]Gڋ
�2g�7�S�z$����o��,-[���}���9Ο��*����3�0���y�}��;��-{��
ֆ�j�I�ȗ����-$V����w��$�,��T�?��)΍\>��W���|����_���94�g�p��˧ϖ����o�.on���T�J�4�)m��D��e	�Fk0����z��(�H�)R���+׮���p��E�2g}c�(�h7��tp=�0j�e	��QV)���|�uM��2GY�u��(�|[�`��%�F��P(����G�H�nE	C��R9h��rQ�ñ}��UV��U�=u���]�̢�*)���1EU��e�Ӟl��~�յ5^;y���Q(X�prÅ˛l�vuי��a׭�S9N�����u�pZ-�vx�)���q�6X�R�
:��H�r��_fx}�k�WYƔs�B�-��FdЀ4�n8]r��Ont����
NQ`U#��/�N ���&uk���,B?�4��2�?��&n�v�eiBVh\/��S\$�u��da����9���޷�����~���E>�>ϯ͑�wcZ����︇�>�k���Gx죫L��[�''9w}��x������~c�2�� gW�ť+'�s���Cǀ&�=v�w��|�R�����V�y��,?��������Ͼ����/1uǷs��Z6X�P� ��@�C6�QV9:� /0���U�v-B���u���4��Ko�?��y��
�^��/7;�W7Yz������v����R.�QF�䘲�;�đG	�"�c��m��l%	\�FvX�BU���u.������Da�<�aH�xTF�l�����`T��(t�(s]����!�%�[�]K`�BDUQi�1�V�ϱ�-˪�L��@�1�5QI��!,�&j6h�>���l�.S�R��d��f4p��5��\#�S�(�hC<�1=9��v3���\�xًI�g/��No��'���'� /��A{7j�6Z��	�f+l�6x����k�q�B(Z��	�l�[.�Vl_]���%Μz�z�6��q���Q�=�����qZ��ph�VY1��eО��Dc
*C�+Ja�������0��Cl���"��|�@'��`mgi o�6S�6X�YJ8�&�oq}����~��~`�ç�r�?|z�gF>������~����O�֟���z��»����C�>���evH������l@���F0�h7m._=���i��ڋl?�����5~�O���?q�=��߾^�;���/��O�}����]<����W�4�6�Rd Jl�B�R9YV���0Ii1p��[3��_��羹��3���i����J�������#z�� �*I�n���,�4�ix��`�u��T)y��%)�4����<�����������p}���iv-���� ,��'���pH�dX���n��O�QT�4I��AZ��_���H*��@gh�՛#%A�c{
ǒ�%(�Q�X����T:õ$ҭ]�H�1�S�G�f��yL�'�yB��yBQ(K�!%�����cvf�0l dM���?�c��������[���{���;�u�a�c�dYʾ���_��-*��hO��7�o���M��$v�@���7#�F������+�9����<��d�qBR���s(���*1��j���k�A��4�KJ�6���@oPX�qAHl�ƻ�	qv���A������]c��83���[ny(3]'�-�$�a�I�"���W���h�`����\���_�穯G��Cp�1���؛���eڍ	�������d=���u?S)<e1���d���g^�iJv?x+s�����7C��	���G�����}������W����ɒ���]�q���
���B`C��s�3~�������s�>7�Jt��G���}8� ������u�X�ڤ���D����dH&Z-,6���S�؂G�q��^����ͷ��������Η�z��˫��$�����;q���k8�K�ٔE��K�H���6�a�q^����|LYRU���0����bw@h�M����[ʪ �t���)R�f�x<���5� `cg�,#��b��R9��TT�2E8�lq��!x�N�|�QdER��%���,..�E.]����eU�??���o�6����铼��+l��T�"�����������7�RH�u1R!,������xQ�Ng��Bu|�R�4�k�s���z�������H4�eS���k- �(����*�Fd#��[
�O1ݼ�r�"��&a+��,!(}Ӱq3���3������b=mӞYdu�:�SS��0�	�ʁ\161.��U�-+g/q���8���sםL�3wO���4��:î�\�~��z�	m���m�YI��T�H�(r��I��%�gx�e����M��U�p���a�P�]��f��9~�^NY"�*�~������.���5�R2�	h����+�ʟ��d��1¡���r�^}�O�?~��,OW�O���_[#��������E�l���BX�2�0���iU1���XU�MA��q)ٻo7�벾����
�n���~�#�������g>K�7 �KҤ`kg�$Sd)��m.�;�{�����o����m*,J�%i�M9 ���w��L�[�>�S|�7����X�d<��CF�1hM�hS��)i�p��)�͈��?ί��/1�mմ|W#T��**C�뜩�Zl��?�C��_��_���/�%1q�P�q2&�.]����uF��$+J����+�����z�I*І�q)l�k;�I��h��ƃYYwV�|��Q��Q?l"����#l4�݈0r�KTN�௯��Y�l��&M$j�2�S�
|��m;!��
iJLep����3/ъ���b�!��t3�b�$�fZ�t��UcwIe	<�R��,�����Z>+Wα��6�6TZc6��!�H�u}v�FZ�YZ9��!K����9��6.p{b[!�9��*��:z8�*��������JW5m�`av/��<n�`y>�LQ"A���<�ѐgU�#wolӻ:b��e.��Dw'e*\�S�[C�t��ZKDe�݄[n�?v?�xTU�y����c�)��X��6X�\���f<���MSg8J���YpC\�����C*n�4S_ap��,�%,���]��A���A������a����4ʲȳ��,�n���nwѺ`nn���9,�r$J�o�8M0��,+�2�(2,	�Ϝcaq���ifg��#&&:�F'���O��P��͝\�f�x��{	����H*�<�(r���	�u��?�1�f��N����ɩ�'�*C��Fq�B�PT%�v-�q��'�$/5ya8r�����n���*���1t�����S��llwپ|yC5h95�L(��zHia9.��k��t��(�qu���k���pq��ݷ��W/am_�X dM����D�
�DW��q6��`M�����6���x��ٿ4���B`v���>Z��`z�C��y��'i��af�37MZ�,Cz�<�����ώP^D��85X*���iN�3a7c���У�D�$v6&m���G:�I�1y��+C!��In��^��f���'��J�0b���!����<���񔁢���StZS4�2�p#E&6{��(%-%�$�|�g��~��م#�;��{;��d���$��,�\����V�+�F�hD��LN�a�r��o���$B��0EN��)M�������'*m�����'�|�q?�[Ո���M~���-�?�O~�iF�P�i�x4&�+���eIws?rq���E��Ƕ��l���f8bY.�����d}u�C��:U^���@5���QdE^�t%�-��@�U��N����+\<��$�����6�*UVҊ�����/�����qB6ql�4��a����>�$�1+��~�Y���O����}�Qj�h�#����GN���7��vm�]Y��]����J�86��궓R %�q�lۮ��B:�v϶ټt��������6W׮ /_E_��5�$M�,C�
�s?�o?hW%��ST������;v��{Q�Ga4w�8���gYO���v�E�gx⦇c5)ʔ�������p�k���?�V��9{�'���g�Z5��嫮&��I�6�rA�S���w-2kDb�7G���v���ܣ_�����؃D@Vr'"Q�P�J��0��N�@$eEј�P)��%)���[�����%�>���������u�r�lɈ��,�s�ܒ\d�VY����$VΨ�g�6��&���G�"�ǒ��(��2�B��y�@�e�7�iF"�\� +zVy�߽��|���
��5�����^v{�l��85Ao{��~����;L�p�i�g%�q���$�dD^U4"ױA�<�y�'�zu�r��8NH�(�a0�i�i�򔊒�����?�?|�Kd��q��9���ŏZtG1Q��z�6��;<��'x�+_��S'��� �J���RR4��.M/�����%#��կ�w�i��������A����eY��"4��={��zmK*l�crf���Bc�r���ogs�ɡ��lm��e}��}��¯�$����9��u���.T�U^0��Hu�-������{nㅁ��E�I�7aH��{�����$�oxr�D��0�����?#��l�q�t	�C�O����
o:1å��/��)�h�o�M(��)NW�Y27�aomp��^~�U��-<���g[,>���t���w�Ϗ����o�k���5fI������l0_N2�,�FP�	"H%l�=��0Z�6U%�(����$��h�̲)Px8�h
�,�P��1%p2pD�TV�3�#,?@�E�b�ےS�ܰSUB1��e��iiJY���RҴ$iFa�r�4!�DQ�X����*�4���i(��Lpl)����+]
�c]笖�K������s�˴ϼ��Ľt�pZ��H�V@���e{{�5f{+�((<Msn?��V-hz�c��xiW,�Sx����XkT�R_8{�%�a��Vs�Y�;C�4#)E�V�;�RX�&+kP�b��[;9Ӎ&����!&�±�ٳ�e��Ω�wc�=��L�e��t�2یˊ�m���&R6iN���5Y���I���oŝnr��.]<CT:��ai�.R�`�p����s|��Iy�9~����&���g��;�������m?����ŸB�n5�;X!M�v��/���/p��y��C����������ҙ+8�ԓt?�[t֠5�3���߀G�]C����g1/�H��~F2�Q
;{�ĩl�ŝ5�컙��+�x�h�I��*b|K��[��C�>�u^��Wy�̝o���K�D����̍�l?�ы'�T�L��FN4-ڰ�eqԳ�E��c͊=�Òo3�
�\�9�Y�Kvy0ߴY]�<�ݎ�\�b֯�%�n����+&A�L�%�NEǫ舄)�2k�L��)�dR��
�����4�nEǩXnx�1D��W�	G0%rf��iS�˒�+	���2��h"��iU�дeE�*��!*ƴE�dP�#�VB(5��𥦥r����M=�'4U�C��b:� ���*ű���)7hw��^[�Z�C՞���&�rH���C��J�q�`c�T����v��u`0@�CFF��a(k_K�#�N��d���C&��[�ݎMS����llv�9YoL?OU�� OY��=���/͸VV����4fk�i���Ϩ/��v�̈(�1�3@tw�=����ȼA$}�qL��R��0���#��N3edI��JLQp�ޣL{t�1�|�Vo/���d����\����d�o�<���>vR�ӯ_Û��g�������X~��m_a;���
�^{���~�6�����y��7�-�g���������e�,��z������~����P0>��s_�%# ���I��������f��>�Q��ٿ��/0��$�h�������X}�y�?�I�h/������f�f?eםG�,Dgϰ��O����Գ�:��Z&'�p���q�!́��[�R�Q"�c�,�/2����pr��9�P=����F�e���RT;ECSl���{X�B����gC���*��NƸ�a��(���,�.&7(e(����)�d� 1�X��"�����Y��*7X���)���x�V��R�U�)K��@�<+ɪ��U#��Ū�I�LJt))�d�������Ok������c�'��˺#qゆ���=2c�.���h�P�HMe�,.�a�*AR��j;t�V ��j(�_Jv�����Á�D%��8\�iL�<? �q�e���Sn�F8w��˫�<&��X/��LG�/�4C���c,Rc#��5f����M&�>�����za���x�2��LRj����L|��[sZ���Kt�@�3s���
;������p���:�(6��x�M����7p���Z�˞#�P�'��cO���ؿ� �?��دѻ~���������.1�r���7^��⣬�����ྷ���}3�nP�����W�Ӗ�$	a$s�;�?�����-`����������k��-,1���l�Nc�m$sGt���7؅63��_�,���������o�f��2�\�C�ϼȩ?�3��m4~k���=��O���a�rIU��4����]),aS�5Q\JI%+�T-��*��5~f!r%�h"M�D�L��W�l�6)s��c�E��OaB"�`DVD�G��]�
�2�2�le�������/��ad
W��H(�����"59i5��4E6�(#T�b
˄�®]Bn��F�V1�\3a,�SI�J��xňNr���<�N��uf�͵˧I���[�+���� �\<ͨ%9��Le}�|L��_'�m3UeL���b�d���	t��W,�6G]���"�;��6��6�x�����	U&��cv��K6��-,���f�	�b��LY��Y�$��1{�fF���O�F	J@Ӹt���Ϥ�҉Z�͒G��7�6zC&$4�!b<��4ƌ�'J��eʵ<01���]ei����:�/s����/}��tG��-^	��,_:s���yy�s�#?�ɵm��\���:��I_�U,p�u��Vq1k![m��w��inYY��W���T�AO�X;%�`���߁�w�t7��a�o~��O~�<�p���4��^ɱ4��6���/�bvv���6����O�D����Eo��W�g�=�Mo��r9�j�^<ɹ�֩KL5��C)r6�y.|��sf��l��F%���)����'IŘ䦢��-K"��s����C����<ec�������Ѩ�D��=��KM)m��J �$�K\2�E��hD�$Fj�<&�$�2,m�ݠ0�8�¥DT#��,*�J�-E�K
K�R02������ؖ�������+�R�A��`�8�)l<-��"5	�(�6M3bO�v]z��Ǟd��t�xWW7JE�ٔ2'NFl�:���h�c��U�'�<Z���\$����`�s�r�w��F���c�U�l@�zv���Qz.FؕG^V��%�M9^�6)JCYJ�T~��r)��_e�&�,2+�#J�x���r	c�Emz�Kh+�,E�6��%����(�`�����}���-P`[.�0;鱽�B�!��hv�ũ&snIZt�y����O�$��}�a�]�pￏ��c��s�$�}�[����}�x��d}���Q�Tq��0�����	~{�e��=��k���ص� )И�k)���o}���4V	ݏ�	��4Uӥg4r�Q���lF����{ӛ�O���1I4G��~�1��g>���n���56����7�;�8)�/|����K{0�Ӑl���q ���!�Yz/�>m-�Ԑ�ht��d>�T��T:�)*�UJ�Ht���%ٴ���0ia����h��%�Գ��
2��V%@WNNˌi�=ڃ�6X6x�Ms�M�u����X40F �[��̈���J��-��ĥfLA)
n=����.a�)vX!��R5U 	FJ�?&;d=w��n�<���
�!'�G2)m|e����{���}���#̞��A%�s�0��Y��J�},�%���9�dzY$�yNV�L�q���\V�����n"�y"5�űʣ�i(C����;jQ�.���l̼n��)��ME��aG�2Ò�d����خ 10-R*rK��)&�]���(
��S�&'g��7mi+��F��Bp�7DX��!��,��x�)VVs��|����{q�Sҝ;�(��e*eTl����cOp��9�M��n�o;���}<�Э,�'MQ��#Wqn�*��۵����r��rK�e���1_y���:К�$��Y��o������Qt�M���?���P����A�+�nE�bަ:v'��G����]��R�IƏ�=������3��Ж�S����	s���
$V� ,���~ؾ�?��� ���o��"��%|�T��ʑ�E������U�<�-��9*�3w��-l/"Ir��jM��Ҡty�+�T��MW
2i�6"7H$���=����c�F�d�<�<�ȃ����T٘�#A�(��4�2-@*�"b���=�whx.V�Mj$x�8n=mb{��aY���B�Js�ܫ�[p��
r��3Z�,�h��o}��+g��L��000{�nnz�m<�ͯ13=��|����0���Or�������*�TX��j����໿��`�g?���-+�;�ⅿ�]�jAX{`k���M'����n�g���g?���Y<q����S����v!��н�m�۷�����?�W��Wy���_���/I��z� �n��<h��tvs�ŗ�l_�����n6?�)�u8��^�y�(��|//~�ܺk_�������A���ˌ#x�7��Z���*��F ��u�!�s���2��)^�_�RXS4�y,�Ed]����8f���ӣq�,��k�]�P���HRK���Qp�kp�g�~7�?��V.�ϽH|�q\���kګ��tW����x�Ef.^妝m�(�u����œL������H��XY��3[�3�0l	Rc0��kS!��7>� _��"/<F۪����K0���1e�<^�L7VN�6�W��� ����]L�5D��X�*bt�`�Q�**_��	i�::���_��^�M�1��9��&�Fɂ�I ��]ə���):S���r�1�2I)=���UV"uE�n��YRg>{]����&��U�W�2ؼ�Ε\z�u��9MUvQ�e�K��%�U����>Xa���Q�!��+���46x�o�R�ye��{�ŏq.�D��c��]��ٗ^�}�X3Ӫ��E=w�{����3����r������#�����i����K�W�S��>t/��7r�w=ʥ*���<��/�}��}�=���n�+�U���[�ڻH��A>p�|���.�0!ٺ�܌��q�0�� �
��G�C�t�6b
��c����l�{�I�� � ���̵��3g����g|��i����u��8-��'_�ui�QT0��OZ`� �ֶ)�_Ļ|���wY���!�Uk<�����&w�nr��U���E�z/���Cd��d�]�iK[���U+ �|7f����\j�~⏉���X�&(�u�#�U}���&I*�DCU�@҆qV7`���C�^p)��������4���0�h" ]��x�>~�7�����.`
���*1��]JYY ��F�t��I��%�����&�R��Ieji,��E��]i\�CZd(�48J��Ԫ��T�6$ʒH%�)�H��j��ض�,3�I�g(c(����҂i����_RhLY���A
�6!�-����AQ��ԠmE.r�|D��2�F�{����8<�1����C���-oy'��'h�M��;���S�z}n~�Cl��_r�S��.�6V�d.l�y�o�/�v��Ɂ���+?�����y�����)��� 6��w{�w������������O��K�92ex铿�A]�����5<#�y����3��׮s�]'�?�����^��Q��&����}�f�[:���2?k����;Nf&3�L�ͤ�f�a�M�X�b�)�U�h�����bE����RЀ�s�jO��BӤ�I�LN3��f���>��;��Y��}��{��wY���x�?s�O�!�Q��Wy�ߧj`ԇ&�y7,<~����4���,�{�;8z���_e��q���x�7������W	U9a��͎� �	�qh
˴�6+:�^:�U'��4� �u����@�t���^׋�����Ǿ�I{��H=$�)뙃
h����8��{�A�K���,���'��p��}K*d�O�
�ŽE%��K)llN�@I�s�p�T9Ȕ]kI�M2����3�1�8aZ�$c��!6	�n�]����3S�%�=�*�H������8�x$uS�BK��V�"�V�EÞZu���TpJv줰u=�E`�}vm��Wnl���:X��Kb�£D��@���W�IPң���[ʶ"�<R*L�$1�ш���C���mj��V�6��aI�Ҩ1���5��#��A�R�S~p��yƯ�,�O��� ?�ٳ��+'���Yv�:2�LXYq���Y���'�|����:G֎r�ԓ7/p;�����(F���L���	�W��J��Ͼ�`�����z�o\��2��Uj���cl�^����͌�~�;N��<_}�AK�ܘ����'�pssT.��g!�\=�27O�q��e���˜~�I�)$Q�7ɐ���x�n,+�s<����;w�c��:�)�t	y���可r����딬�B���t��.pN������ �%�rD�P��ԧM�M{)� c�uӨC��Zj)0F#�l+x5�z������)E$�4~�A�U���x��W2�R��FkT��UЖ,�XJQ��g%�J2m-�Q��FG�^�DT���	�N~�i^9�{b;��^'2%;n�D�!�!oi�ge���l�g�F!�#���U�J{X�=H=��uk�*��-��&�}��LK�mQ[�i��&��Yg� � �BYPu�.
t1m�&�۷���R�)-Ă^���]p��F�b'�e��܋���1Q�2�Ʋ�b�n����B.�0Hm���?�%�֯��Ϳ`{�va���X}�(�/^&�S���M���p�_os𓫬_~�����CE9��W-��V�����{l�s̏�����d�n2�0�c�lBjJ��yF�s��ER�͖�Ճ̏=���5��y�)B��23-ȗf���Y�U0��m�y�h�g��5FT�;T�I��H��}C��ȱY�5]��6��R͂���%�����H�h���GI7&���2�}��$��v��K����Ѱ������>�-��2�٦*r��"!�4q/�;KY삳] ���aJ�T��a�Q����*��c�����b!$�#�i�>������=�    IEND�B`�PK   r��W�ѿ�*� �� /   images/73de3dbc-74d6-4bf3-b63d-33bae631b402.png P@���PNG

   IHDR  �  #   ,���   sRGB ���   gAMA  ���a   	pHYs  �  ��o�d  ��IDATx^����dIv�~����[2��r�̬�Z2����h@ 	��h&��$��4��FO3=�L�y���1�hl�#G$`\A#	�$@�4zߪ���r��-��9�p�#n�/~[�/׺�*ψ_č{}=_?Ǐ���������&m�c�0��~��Y���_7�����A��a!�"�Y�jW�����c�}�������:Da}}y��W�Ƶܼs�A��	������0Y��O?�@X��>�{���=�=Fb�+�7�ȁZC�:�@L�R�:-У���Wr�2����W^~���E�}�6�dŲ��ְ���d�/���7�{R�n��[�w��00 (ٳ���"��]���8�ȯ�o�tp_���3W;q�����%�#H�̉P�>� ��0S��P�5'%����}�+�t����|]�p9���a�����/ �_x�677��c)A(�,�����w��Qu�1y \��n {�حv��n���7��e�GO��7W���Y.����(
w��
���~�r�{�]�[���t �hv�@�@MLU�mP� �0������]�أ��#UUq�ȅ�lcc���mL�X�l�Ȣw����g�ӿ9�^�;A5!E� ��aO���ׁ{�1�n�`f����]X�V�s���+���N��?ΰ0�
4�{����.�����Z�@��u��N,�r��0ӑ��ٵQ�*�*�8���A��|��t&R�?�����UL����Q�|�:}��?����XԾ̏�'!D�_|9�mnl�=��ԈU<���-H���~af��d�ƾ]`b s�	�o���a�� -i�>��r�ei��9?^�n�Z6\����^0 ����"��l�a�u� �FAE��r=O��EBT|Qra� qj�;��-�T�gS�^r0��  `Y�@���lG{hy\�2���#�p����E�^��qF8�{�0#����"���_&��`���~�qۘ�l��@��`	F�{%M�⇸`�ה`�6�~U��q���5�"3�H��.$���i����^矻�����|ٽ��"�%�����?̈�<�&B��4�לmyB�hyAZ�kI9�ݏJHy����A�X��T��=K���G	A|�ꖾB���U�bQ)=�����~��e��=�(	��'��a�b��Z�Z�ZD][��q��=a�����V:�6G{�E�p�:$*��WX���ܲe6���>8�ٺ��?EI(&���4�T�M�Ҫb���B�Ns�%IU����أG�mbj�sg���l��D��d�Y٠���lUv����"�ͳ��j�)ڽ���^�6b����$T�V�i��9oSϋ�I�g6���Mj�|-�[_�:`��z9���� �.W�l?�]�t�����_!Mrv���нroY�!���@���a�|���J?�C��*�!H*Q�{�@4�}�z���(�����S��n��է�[����]~݃�λ�L�;�{��=(��/>�8gm^F��U�i.]��<w�9���`<H�M�{'Ӣ�{�u>9j5q�)���o�݇���$��$i�f���9�5)σ�i$ I ��	�׫���ז�a��4j�~��d�5������aA���2��/��0^�ՅCo+DC^(O�=�I�����bV�Z~p�����(9?(zY�,�B��7@0w�+�7=4q�
mڅ̼>%w�?����x�K����b:	����J������t�գ��#�ښ��7�8��.u�*�f˻g��7�<D����Q�kl.@C��p��+�d]n�&4sm�{U�	�
�i5� �#!c�*)����FW��)8��I{�l��R��lΞ�������-%���2P��ۗ�$�ɋח*�H�y)�W��a.w%?#NC���ڶ�m���6+���5V �u�n;��<�版o�w����k�S��}�o�zN'ゑ��)-��gB��W�R��,%O7�w�M�
3�һG�|�Wo��Ӯk�dI��!T� ��.N��
q�z��%�Ye�}+{/�xt�o����s��y��Q�?w`�q���((i�宰����9�\:`>l�זڎy�G2���ɭt�	f��1*�z�,��/A����"�3��"���RHv����g��l��� fQ�k8,:W��[א��'C;so9Ee��%�Iu-4,��?�� s��E���ç�3���J�$x J��E*���~����� 8y��U�n�8��S�8}��-��5�z�X��%N���QbֽKɥc����A���G�R]U��F�RK�y����q�eU�iZ^}��q�� =���o��&�9ڜ�Kg�u2߬;�ێ���x��fI)�9���p+��W��~� ����̈�E=���df*����~�Q�����u�����B�&X'_�nR�Ե(��r �$�d@@PZb^��^�˿�5�6�K����0�&	K���Y�%B<cޗԭ1k��;Ů�f�ߥ����>ح�ҟ�8K������ ��--e*c��"XH��^�b��}��`�����hh�c��b��^R���T��Y�g��<0̬�1�>����iɱ^%fS-n�.���Tey�z403ڦ��ES�q>��4�Bj�FLn� �8r����aB^�ݍX�n��)�
⚂��=��m��n<JH�9��[>[ f�23����M��f���n(W��^��N�3��s:d��Bt}˂�H�u}m���rnq�������Re*p�9p5#�L����M��5�4���O�gD(�ki=�WgN���}#eg6ˍ��y�;z�܅ h00wj�%��+B����cΔ�g��gO���ӛ��1y�	ɟ0]0�tfZ�.
X�ҝ��|��'"�û�w��g���e
	�v{t(#V�2`�������;_++�Q���@M�I���q.3����%[4��|�yY*-&F8~|��`@����!ìSI6�^��.|�gѴ�zPL;�5yq*[�1w76��ܜ�mt4.b]qd&x<;	I��!���J��#U�!�������4z��o�g���ǲϖA��+�ٿ������I�6$5��%�¦P�b�7R�f������f��	�t��f2����"�����fP�51���2�*Ys^�S;+ĵǽ��-
��q��+}��hS�i��c��	M۸�[H(5 *��S|���[$���ҝ�+-��"�����
1��k���ш��&�8�Ɲ�T��!�ׁ��/�t{t�.^�^�`�-4B��?b�ж��d�i<f<n���zڗ����uj�y0�y�Da�$^������!y��8x
�E�=�\��j�kCVW����:u�Օb�5U�Є�i�[/3��O�~�Y(I&�Z`�+��.���0u�j�nlr��m�߸���&[�c&��Y��M�dp�@A��Q�!�R��5QEX_�9vl�c�VYj����V5���!�^n�R2�	���5��t��s��,��k���G�1o
��B���7���b{{��;7���5��:��s������NJH(c5JMKEM��ňւ4�����r��1�WW���jY���m��%�]KrɖS�|m�53��R�.$�K���_��6ܔܴ[�mnݼ�͛7�}g�퉛��"F�M�Y�'a⫙�-�f��� ^��m�1`P	�k#N_���c����2Za0���)��.q���{u��⟷���|Q�h�"��`��������[�ڶekk���M�llq��w�n��ݠ
F����D��d��ͱ;{�h'-�^Yt�G�t��B�G�D�`��h#+x��K�������=y��U���uf��	d3�}�jv��c��^��lR��˰�Z`�$nܸ�ǟ|�k���{�ǧ�6�-����
�=c�N����a-�
��Z�mƤ������'�r����'Oce4p�p� �(�`��Rzŉ�*�<�"v鵋0%?:��W�D�� �I�9�N�Ο,$5nݼɭ[����5~�����W����4 _?T�N��kb2�H�!���H$����ml�.=˕+�p���8yb��ʀA]3F��=�URRb�9�o[�!�eI���g�na� c�T�.PM�*��?����z�����w޹�ֶ�oR�P�T�R�DB|�w1���iAdb�B�*�lh��Ǉ|�����Ο��p0dmm���|N-!��r`��1�!��P�O�v������cw|�X�`�8��h'���-�߼�~~���)w6`<�~8�����L������'Z�m;��3������'T����%M�:w���r�Y�=c>�o��������9�����r�"_<�h2E	�)m;!d�B���w�E!���ch�B��jA��R�y�MbFV��b<V66���k���[o�ƛ���׹{Z$Tuv�w��2�B�&a�a�n�6�y���˯���+�r�^�x�����D!*�"��ݒ��*��Y���eS����Z�]u�f�9c��#h A��Uq�w%p�Tܭ}<i�ܸ����ٛo��o�ƛ����-�nVl�U]�@��g�� `�Xp�D��0���i���V�/�����r�E^y�y����6�
b45���E;=4!��Qa��e�Y}�Rw���t�nlq��R������x�h-�ׯ^�Ï>�wn����;�������ꚪ�����At�q}�18�A��`�4FUms�Ā/��W���+�x�YΞ9��2�����6����"���7úkU���?%w�c?x,k�1�T�-y�n2�a��1�#���
�%FRRn����W��O���7>��7��杖�8!R�Z� �R�����W<b1��a2ix��Wf�9��&�꞉s�����;�a��+�n1�`
�p��:��|�������������p�쳘m#A	f�&Zi�W�:����,��aG�XBB��[Ԛe**��h�)f�6nt�n�a�x���x�g?�?}�o}�|�����Nfì�4/֚�Ex���8��q^|����/��s<��OgTMj�f�ߢ�#��Ȉ�������B�?��K��0���2A�5�k�m4�d���Vs�	���#��17o��ӫ����^�?���|�M>�t�ݭ-b]c��kKr�Lۿ��JE�"�M�6�<����N������r�/\���Ӭ"R���Xl�k`�^�����R�`�G� YX�O�Y�g��wm�D����u�:|x�������7���op��Eb=$��ԭH�P[�Q�l�@�b�#��aeE�r�_�����_�����>3���4[��^S5$b�.SBgL.��m�/�3s����tH���x�ǽȑ���<��)�aM��A ��ֶ���[���G���w����!�}x��7�Ҵ�
5đO�MI!�>�W��}u?�<�I˫���!����(�׃'Nw�0QD��޻n]�'�"����?Ǘ�t�o��/r��	V�jh6�T�	�cʦ��3�Q3'�ˆ]��'�|J(&���%��\��ń�0����m\��e���*R�\��	?y�C�ٿ�C~���\��H
�#w~ك8��rNR��-'NT\�t���������p�8MS�	�٨Du���a�&�i�m��+wG|�d�^��{I7��0�7L"1)*��@
F��66��f;�my����:)A�cVVV�������>����?፷�q��m�*,��줋?_\M�y���5�-��\~�������o~���3YU�4�Di�0m��*�2�@�6%����(T����eR�],�Y���-�?�{?�{��ՠfe8"h�pgC�zu�?�������������Yի$�\�>����!������x8�y��:���/�.�te��AK#&����b�����[�b�5�,�iZ,A�-))枒��P���
+y��ѯ����̌(,áa�*mS�$��?���ѷ������|̭[J
�:�B,��"�:�������APQ�8q���������7�M뛷L�`E�Y��q��	QA�;{�����B4$�}�/�/�t��V�n�0F�a�(�*(%��H� F|W_�KU� F�1*1��y Ps/^Q�@���9�(��(~�F�	�&�l�(+� 	�I�M�� �12��'-�nݢM�f0]��Ռt��u�8�)��x��
�^y���W~���O3Z�� Q��B/��f�FAф&@ʂ~����h���K3���Q�Pk	�"�d9%wSE�E-[��D��-�;���j)k�ZC�l1iZF����
�nor��6ׯ�¢�2 H1��L7˺� L����d� gN�s��E��s/s��N���6��Q�6Ĥ�k����4n�)k�|���jj����?T�v���fE�3J���yW�K��[L�U,M0�����l�����Ƅ&mR���ה�pߜӱ�,�T�2�ѹZ�}�8/]<�׿�s\|�$ǎ��*[����'1�	��1�u9���OՈfTfH��Y�O<��m@�C����Q��Ѥ*�Q�($"��h��F'yT �C�_���;lnN|�X���h��wX��z����:u�;[[szt()@�6��Y�d2��|f��♓�?��Osl�f]����:;TFq���(/1V�P��Xa�0�v'�(�A��V�B��w�{��54�"�k�U���fH�U��Uڱ�N"U��y��^����_`mmD��%�r-���HJ�@]U<{�$Ο��K/2ZRʎ��M�����H����������71��1������r�,��%�1����5A�w�5�����B0!d��T�U��g<!��Pk�Ξ9��/����u�<xE��HF?�[�;���
�#�9s��ϟ��/rbm�'Xj�&499Y�`B*�@
��")m6��\3%E%�H2'S�Uɦ]�����D�D=��BB|�aj��IT���u���f[i[�i,��>���'����:}���P�)�rNT��yP(uϞ\���3<w�Y���Q�:4Ar�l�7��(Ym��<���7�hyա�L�D�t(g�)K�����<��N�n�l)�0�MM
XR,%V�G\���=˳ϬPE����~B�m����w5(X�W=���	���*��!x|˔L�g�Y�_��O� V���6�� Ê�	M;!��4m�X�R���	����[3H����":q�ImJ�*)�ԯ�A� �Hڀ&$5�*��TaDlk�Fi�ê&iK-���8{�,�N>���*U,Ƭb2��k��a�������8��3Dk1�r�\ۺCH�����*,@j,Z�*�x����#Rb�8 ���#x1U� �\�a��C�U`(���(FVCd���ud���԰:�Y�k���M6�v��0p���N��̉U]�y<�-?1df�!�cǀjPW��ϝ����1i|��x��Q�@%"e�R�A5!V5� �:��2���I����іFmHڐ&M�ȯ���䗒��sc��x�I9&��v�PEB]ˍ��*e�勧���.��s����	a�)����1���8{�$/�t��֨cKj&�N0�A�\H�1*�=Ւ}���$I���z�=�o)�Y`^�m}TN�FXr4�n	���d�x��V�Q&�X+bԡB�Pa<w�gO��g֩k��`.?MR�q{+R����@�($f�nB���\��ޱ�FCN�Xg}}�����A�p�(�t�D�Jmn&D��r�E�-��C�v��N��$I3��3k&�$�4uH����Iɷ7����?��QK���èB$Ɗ��Y*���jC�I.�R����Ο��/��a.���`g��=�ݑn[RaP�e�U^5��z�T�j��;��c`FmFmBm���&�Ja(Ik�Օ:ek�����@а�84�S	����:dm4�b:&0A��{V�D�<�+�%m�Y+�
��ި����BI5j4־-$T�\!b!B>���"z@���dq$Q��E�����RW?�
!	�����Q����Օu��7kI�s%�ɫt�L�GV�����F����i$c"�3�UI�"�Iu�>���A��1�'�l����N<@
ɟW��eJ�*x����v�Fƃ�rx�g)�lis�J���B��qa���6>�=�6��ԕO��������=87���uf؏
��<P�k�N�8�y�X��pX������*�����ZN��ͽTS@%��.�h�V��׸�C2o΍K�o����kDL\��W�tŜ�|ZGNR�ɂ64!6 JJ-Ե۠���#��r��3�&�*�L��u"�-�z�P���rǵ,��ͫ�`y����KrB]��ƾ���I�n7�&3�D�Vm
~֓7#K��'4'�j&�Ե1DZ���fr���lOp��I �u6���V�A+��n�4��u�
Ai���+�H��2��C"�WKD�Y��ͮ�q+F_���]e��:��^���1#���u�>I�A�WF5�a��\m9f�o�*�t�~�L�!
u�5U����6 Z� �j�a&ШXP��z�=��Ĕ&������J
Hѝ�ڼ�
��e���|�ނs��'YPBpӷ��~��O�S�|_-w��>5�R�:���j莪����� 矼��{���\��h+g&8����YYPW�%ds��y�(��\�F@S��w	y�0��n$�Y�����S�+gMT٥M���ƨ3��@����IIR��T�M����� �|� M1��4|Sq�"��e��ͤqGq穐g��aK^�C�y�ƒѼ��0E��/3���V$�"	�XpG��-!������F�{�%ѶJ�
mm�ٳ��L'�0����Qh��G��<�>�(�A'�TCVG�X
�F*�1���)��Ԓ3�$�К"��B�N��-��MݒВ�%y�r����G}r�A|��	����@U��!�z�vQj= ����-bm�H�@h���`�Y{�j߭3�p�g�m�6����CM�FED�]�@��gkB2��R^�N�4[����QNŷ@m61�뿐ט%�y��d<臔{���ه���IM<x�g6�.c[[1�g�lM�6��c��E�vIg~�(=z�0��Af�T�Ȑ��B63u۹� 7ͳ���!%d��ay�{5���R�}�-IQ,ż^RX��󏂥ljN����VQ���E)_N�hsfj�=8!e��R�S2(��ĩ-w��򶙀��m%�92w�Q!M��"������g��ϗ]R7]Ɛ#�F�4J�k|��S�J&YO��I2Y���!���:CѨt�<��S3�:#�z������ �����r
yj޻X��+�-M���̙�=�&�Xַ�Z7�����"�L�	K)?ӷBYJXH�$X1G/����{�fzR���?SM�m���������H>4w�(�AU�z�0����d`YSk;ڠH�RP4�4���m�H�?��dW6ז,���'ŇoN>�rO�å��YJ�S	B�U�L�Q�Zz�F�Py'1�䱩}��(;1�e�c�F��Z��6:�D�z�Z^t�*U]@������7o8���������B�C��ea�t�$�����M��}!���\h�% �����r�AK����+j��
	�(�U�p��d��'~�S�uUOOA)d�J���"�=,e������7%�$esVr:ydG��kIm&�17��FS����g�!z䐙��8"%��d>M�AVAjbtOj7��9���}נ�IZ�5��M��b�P� M��������%�ϛ�HLFL�e{��f�A��d�Ը.V�2A�͕��ֵpk1M�LW�c�9/pJ�z�,�ۨ�I����y��d���W�� B��(䣤��z��6�䟪<AsV��Cw*�-�O�T�I�P]n{M���"����0.����웰ʒE��M��~�i�T����#�e�<3�g�F��0�$��M��nhq��e��ǌ8�`��y�7"e���RrL+��Xʠ<L\Y��V���0B�B]�Z�iPWj�1�0��0��F[��q��Y�y-��0Dh�<��t�� ~:�dAd>�u!���yg���9�E#0�pX!���r���0��@-J���	d��x��d�8%��`�Шe�Q߷5�������6ٌ9A��R��ҽP�|�((!�3瘅dQ|��#�!"P�O>>��<Q˵25d�'�`Ӊf��b �;����C6�[@��	5�����)m�H�w !��H#!V�Z�*��8V�#FU�'(�'rЊ�e�F9U�͵������y�E�"c7��ٸ<J���_R��n�舞r�L>,��B�����F(1�T�����hBS�$�3<�&$|s�PRR�&R�m�;ù��OH~�C��e+ZU	1��1h����7nr��-��r��|C����K��ǌ8)�B��?�h��s�+L�~
�#sgV.��7Ӂ\4*נ&��m&��	�f�I�ɤ٢i��o�=M[l��N���=&5-���0�5��o5��������F�>G\_	�<[�j����U�|�A� )�����D)�k8�M��\���Ό ds__��!�r�	�*Q����
Õ���qA*�s������o�D�嚦D��w���ǆ�T�)�	9?���\�emY��(cFj�,��u����{׸�g�\��#O��c!#����O�������!؁H��
u]�%���)f۠y���*R;�i<YjA͏��*RI�Z���3IŎ�JԼ�Q^�V�J5�nv���\������o��&����"�[�Ŭ�5�D��$���lbjB�Ju�N�LZ�qz��/))VH�����;�nvE=ʙ����6m3f(��0�N���;����|z�M�1��ȃ�1��F�CGGx�Hݫ���5)7	9����=˚c�������l6Ϥ�rR�����)D|v��𸢚#�4�P���J��U|OX�O/���(�-U�,l-�	�D	��g���̧#��8:q��;͘�p7�\;��*�b�����*��2@�� d��!�D?��*���A��a��C� �~�IB��Ry���&Ypg"/eyu2u�$�qF�XgY�|ʄ%�ɳ� y�H6�R)�N�=�=	3#F���b���;C��h�ř�т�`@�1�q#m��dFg�(�{x�2��d�+1��|��&�*x��r�����:M��᠖O���y-��C��s"����D�s��"D"I*��(��DZ�	�i��mҧ�Sq�����P��!����;�c>�v������17oo2I~*���'?�軏�	�| ���LǮ�If�E�i�`�̐ ��UV��^9���1VW���~�ckϰr|��c�;�ʱUV��uҪ~|���u�`�`8��pl�8+��<^h�A�Y��V�L�0���@L��b���9�Ӓv^ǰօ�L{C�M��U!��sI�Z=n�,�0/���ě4{D6ФD;��>�u=$VՀ�p�`0b0(g|�ً��`��C��*�`�j�}-.�
A��ǩe����R�߳�b�ޖ��:�k�Ϳ'fn���?���!)+1�2�N�S�bʞ��!�q=�D�0�:B�
T�������:k�V�cuu��^!�b}P�vL3q����/F/���-HS���+m^z�Ajo�/{�u�sg��&A9&lf����h�p8d��ʠZ��Հ�Q�+H	uM]�T�MuM]��u>.'�j��a��9����z8�^Ye�����	�k�LRཏ>姯�����G|�ɧ��,���A0k�����s�����lmoQ��ݮ�������Ay���%�sYӛ]�=^Ճj�������U����x����	H�q&-����ׂ�쭙7ԧ���E�u6�*m;���7�B�����s�E��$�EԅiU�0QT]S�L���v]֝"4x�U�a�j�$W�o�����������_m	uMk��i���zY0H��2Z��ɚ��_��_��׾��-*�E|�>�oG0Q߸�&���oH-4��wN��a�B�ڝ�dm,�\@�-	d��,E����森y;:�.�GՄ:*��Λo�7��|�/��޹��-�֨+?�Bv3�՛�4dRN�g�U��_������+��ܹ�.��&����`3Z3R�o7���<Q�6��ВR�i[��EB��
�� ѭ(�"h��z�+_�H<srm�LZE4��'�jٸ2�?�M�=�	����u὏�����?��Oy��k�,	�dG;����4��	jc���_��_�?��_�����&�a��	�*y�^�2�K��	SD�&D��}.��k��֢e��0PW�3`�s��}�g�'e���ack��;[|�?ⵟ����|���w�z�	1"R��$\�CL��C�����c9Yb�4�z���A��\����.����"�&�Z_�
)G	٣0��x�h!j*�צU�z�c67}q�X��p/J�;������w�s�qqAY[Y����������JC�<hx���*���{XA\=�����wȿ�����}�O��H�grZ�7�����Y�3�2\���N�_���^��mH]�L��$�lv�h���
I��Ƙ�w��sw���C����\:]����R�-�7N�Q���ǎ�s|}�8�4���<���x�D�	k���'|�[?�O��C~��'������8�+|㗿��k�L���>	kw'ىM���*�ڍ�ܸv����)��q�PF�{G�����YC
�N�4f0��y��H�6�H�j��Պ�6���o��o���^�N��	��ЈP�~4���¨Uc5��X�������k_���s�F[�8�}�ӷ�y]
��w�np������2I�[u��R�O�\v>%���>_v7Ӟ>�,�|U 3a��&7o������ڛ����ܹc�]\g�s@���'��Q:��35G�W/�į��W��/\�珳2��M���}A�g=0u"Tp�O`8r��M>�t�����zu�v�Po��I�@}�;�솜K����gO��s�y��E.�{�� z�;�k��M�]�8sI���'��f�i��1�q[��;��7��ͷ�c{�a���U5�ǪQ�د�n,z+Z�ٓǸ|�E���W�j#�6kk��cf��A�"cB5PR{���|�?�֏�8��~�o���y�}F�R�#�[/saK�S���4I�˿���ޏi�HJ��_g3���	Y��ͼ0&��MN[������_�E����:��Jr�|xU���޿��S^���ʈ �0!Pc����3��0Jj��3q�� �MU������������7?�ms�_	����*�;�0������`�i�))�Ʉ�w�r��u>��[[д�
a�5��@>i?.�'�=q���_�ϯ1TX���^��$G�qSj�&�r�8q�����6������߾����BkB9`q�8]���iC�D���O��Ͻ�W��E^z�y�ׄ�A�m�\�K��^8h6;��~Ne��1>���w��#����,�ڥ���4��,��h��]$y��ĩ�Db	3_"ִM�?z��~�G|�{?bsK��.�C�!Dߋ7��ݔyo'n.5�������/}��|��V+�4$�0��L�~/����dBU�$;��?��?��3q^���8}k�~�i�8�^��+|��_��w�B��&�Pb�7l/'΀U��������џ���Mn�I�i�V�8����q��H��#(ل���̳'���^�~��8sj���6�؟8%&&M������g�ő��:�Y������%N_^�Т����	�������Ο�����2��AJt'�¸א\�%E�¼gX^���35v���x{���6��c߲��꼾T�
�!}B��Ĺ+���8�a4j�sW^���W��/^������J́ʻ��U�G�XBC��p���y���{�����}6�< �Ry�;׸;���</5<�h��O�/^�W��W�ܫ9���ޤ7Ĩ�Q^�Th��%��uƪ�T��\��ŷ��8�k_��m�I�� �O��A��Qm,b�b ����_~�?�������ܾ��1C��g�L���U��y�DV_����K_�2��K_fm�"�H�:�Puq�!�4�E��5��ni�8?{�#���8߽ʍ�@0�Lv����i��~�7���������7ߧ���a�&?;R��	�E_��=YL���k76���G���}mޙ�*��ٵ�K����{ih�_<������\�p�a��v�h�NT�gP�[j�c�|js�Y!����#%΄ڐ���|��?�Ͽ�c����^mؚ��ҊCp��Z6(o������!�m0C����6�/����o�ݾz/��D�,�5�\�9���|M���0�I�4�2i`c6��;�7&ll�ll'��¸4)�j�K����'�=ΧdX���ޚm��c�$��Z"ysK&�B3��g�r��7�����~�0aq�vk�51z��u����ư5V�����������׍mec�ln�[���cccK��������͠��&��d��Y��?%M��MeK��\�����ῶl���HSv�"`&�w�͹3!�H�Ƥ��M7�2 i�D+�������v��g{[Mø1ƍ2�@��!��Ht����&�Y��$���ё`�l�$Ie�v�x�mm�z)���.��o�l�$p�J��)y�MZh�H�D�&���%�>�1���W�$�G�4-��G�=����҃FyƲgu>��u��p矹u��f�^,ovL�6GRU�H�Y���&T�BBUC�)|cN��w%P��q�IM�l{⨢DBU��UTR�(2��-��[�B�揸% {���-�L������f�W�L����b���ʍ0�Z�`��G=��%a�T#BA�PRa���5����ԨDTI����*;��~�sh�g�,��l��}>�Xt˛������$�B�e�w�$��S~u/�~Y� �FTq�jp�W��U�)GT�b\%T�ϐ�ѽ�̓ث�b�%��Z�:�;׹w�LV�g����
K8z�B����~����C��H�ykʀ�0����$�2�a�t��2M�����V���G�k�������>z�A����Y�t?[�|��3�?R�U���k��	9��7��.�2s��n���-�W �Q ��$�ڟ���X�h�H�y�`	�Ef��Ѽa���b��:������C���tNOh���.����8׈�S �=��Z�ϛ%bF�k[�ՙY˓M?�+��u"D��_x�Wѷ)��i���*1P�h+!d���J�WL>b2�e�)�-*!�:��A�;ˈ�DQ�<�DBE ����Am^;3*4rߘ~T��}L��Y�����OB�|�t��7�*$#j��,��]��C�����*���G�1���=w�Q14�I!F��B�&k�~�G����{Z��/�f���E�א��&ᦜ��1rx��"��������崰�e�3#~����J�,�;1��#J�#	�Q�G���O��<�o�	K�ǁ�Xy6�D���i�z|��C��ka������②�0L���d�\Y��A9���z9l�/K�t�[&�m2w��/~�Q�0�K���>!���A\�N�'aDf$"f�v jZmr'�'X2T�/5AȢ�7��4)3���ƙO�(3���EL.pw��'OtEY�۔�z֒%BeCeF"��|��}��$��P���4�R�M�)M�LI'������ x�\EΥR_sNA=Ư&4��
���m�zF�U(���ʇ�Wcֶ<P�l�
��]�d���>*9�������[�I#A��MZ�l��eܸwӶ4�1n[�'�f2� ؓĤm7ʸ1�|R��y��Q�(��V71����U���Pust��<l�w�ge����)y�^c��^�9�͓f��d
$�U����ע}<�m2ڔ��-���i<pI�&_����S��}���T�K9��jq��_Б��9��H���=q�����U��6`K��/��j*<�{o����"$\��W�G�)Z�G�4}eT[��u)��^������;����w�;w(V��{�@o�?��xם3s��=37�&'���(�Ae�8b^E�3�AJ����y�Z�~.�³��>�\."4�x�0�� ��,��z�<�)�h�1 ш�ƨ(UL�z��?ct��\n��Q���-���EF}��*t���^%zQ�;AϢ�CT�����J-��u�.G��n�-jl��G�V1��������6�e�ˍ`%���{��[�n�ْ�>�xJ-uTqTA�8�ױpf�Dh���j���� ���܉)������Dc\���&� ���ٽ��~9�-�-�U���V��XQs�2�*��U���ې��7����I�Jl%�)�>�R}3X�Pnj�rЉ��rp�t�$[���v��E_zV%P@�\]�Q��g٩���O�H��u���9�C�gB�h��S�+��۠6��ao=w���%(��B���:6ʿh!eY�E�z6z�b5�>�$U���"_�8H=<ҕ�>��ro�8d�g@G�l����S���D�p�Y����u�͙ɮ�Y��a�
8S��4��*�rs�EDmA� 6l�sx�@]���1���1�p-���)��J|����P��糃˱7�,�ns�G
��ȝ�S˛�Ji��i}���ԅW�M�����&����N���-d���	Q����HR�"C���'	L���"�+w��R��v��͚G)V�I��b
��N��*@L�_��q-/�t��'±t�����c��C���{�P��Av�qi-9K٨�X�����C�1��Y�V���>�� �;�O�E�*��oN��_{yP�	P�)��q��[�ѽ6Y�P���wOp��Tꖇ?��8˕�2�R{֖�T
�FP��Ъ����Fs@r����
��H��dh�hж��eb�����v�4I��]���NR�#S��/�2齦e�z�"���u��#��5�~�F�9��3����G���64�\d�0'��6���[zV+ȕCp��9��Mj8��t�v��'S�k���$>.a\1B�u��zVfK(��u]an��q���C��V�J9j0�]�|1��{��#�n;ZK�/�T��\֟�&/?���pM�LfeO��r�7����&������Ӵ��q�*�A�(j.�Vsr�G+3R�\�(6�=�
���K{y�G0.��hּ��[o�RBw.�����]ݢ��lF�͒���Ei�iLj��=�-w�||�kЂ��_7H�Ǚ��#�����:� �M�A�R�{-�|R�KZ�(�U��i�:!�"/�hg�qוƼ��!ə���FՕSQ_$6ʻ�j�����y�.O a.�ڕvS�jzvR�k�^r�^��n:e�ۏH����_n�����^R�5�O�4��sN{\��눟Nn}~�j);$2��-�FD�hg�)�]�O�/P3<�qK(�������x�T�	:��<�*c���$�r0��r�S��z�y�:},NQ}��C^�3L]J(Tp��g D��
����b�LPs:�=J"���,H�+�KU*��e}�m7kd�\6���ẖ�4R�s@.���}Fvc�e<H��$�(ɋ뷎��쟅?�6D����˗i}{�ഽ-���[���찃@5���q���S@M���j�������P��*\b�\���p��`��d��s��NR$����0���풱�ߘ2ySdp8��ovyO1j(%xBHXk�M��Q��	�n����+-ҹ>>:��\3��$�~�>�>rQw7>��|b�6��Mq�F$�̼f���U��&�$�th���ZWK�R��]���'����bG�}���~��)vK9�͗�-���{p�}���y�lg'�����N$Id�ۻp�;�q�HuX��س�C�B��O�I�TAl��!6�%��[�(�D���΁M6yB������N���_����7A�l����'��Vy���^�z<�]S�SF&a�w��#G��&{E�Ʒ�����u�-�a�5"c��9���뀸�J"I!��0p�(o�o �����Q�hv����	��������6��:�@t���6dG�d~{v7.0�����������G^�+��j���I稉����'����!�	E1'-Q��;�&ԾL,�@"䷁�7_U�v5��b�]*+L]�z���`�Қ@�Hp�f;K`�H"DYP�r��ڣ��Yd��cC^�ίL�~��O��/�s��U1�,���L��L Z�uc�1�)린�]����W)�<!�o���d����Y�������������Ē�:>���?_��/�I���g,O�kn���d���!!9 �w}Y$�듰_Z��T����G>�H":>��tIt�"����l~�Q����:��@��=��<� �b�zV'�3���쟨�bS9tOX��VLc��h"ZO��H��C>&7��2
ZP��~8��,""AtH	�[3P�M	|n��߀�.���.Y�l���9�� :4~�4a�C��ч��S�=Y�&��h�������$�R�I�%����*�|��Q"�d�tDj�B��ه���*!�׶��$qb��5�[���!����7�<V<��.���>H"I�4���x.�� ���A��\Np-�tu�>�R��}�]U�����'=ȺH����t��҉_ 0Nn�L�p{�!�� s�^���YH���^E��W�$�7�ڵ�	�|���kmm�	�;�֐��|`Sf�Qqh��
U���,9�H@��*�$zsA��JM5}�\+�N���0	#��d6�j��h�ϊ}:I�dY��D���*�.�M:Q:�$]i�)0Y0_MTM�>��tDX
]qw(>�:����E9�Ϲ>4Cj�y���14R�SA���#9!�7�p�ٶ	,U�0$>����IU��U�䠆r�C�F9���',���g_�BN��+R6<e6�@�� �6tw*T�.��د�q�P��|��)��M���(O����N����@��ӧ���+�S�.>D|Ԉc���t�!|b�~<�7w���
'�CXF��7����L��f�DH�z��=1P����ؐ���mJ��(�fHW�'"�m�)x[��\HX�$�yLH���j��������u@��>�,���hK��$|���9BT��/�����'��}�_/��r*D<���S���0��E����?����u���,��v��?���4-
T�I>~�	�c�b���
3�qNg����h1Rt�{{o�BQmz���3I�O�F�96G~���,��B�3F�]���}��8�	�r����M��+P?����t�����s���m�jrg�䗆 9��uj���A���QF�ߍ�\,tSO���
:F�;l+�"У�~��sq,!M�*�=Đ�b���A�N{�ED�Q{�"d,Ģ�H�jN#�_���8�p�Q]������|���JS��q<��;<d�T����J��V�R�5���m�%�99�㒻�uuuM9	�Ϳ��Ѭ���H�Ɲ��V|)�A)��k/ ��#2�g�9#��m e���1/>B�@u<����m|���?�<?�����ʦ��3Z[��j����%��4�8�y�����O���'m�m���sv��"Rʘm]m}��.1�6��@;�A��$:�������	������n��m�y��g����n�w�߉�g�L9�>O�	� Ahg���~B����"qR�(����f9�
>]���z/;uP������y~߾��n�?������/�G"�s���m�:��}&x��9��X&}�|�|���w��O��g��Z�l.p^n��&F�B�4�߹�K)�$�A�4D�ytԩV��n�_�oW�	����G�s���,|Ě���Khn��:U����������#���{�/� mP�{�{�\ �����3���Wؖ�q�ct�9t���~M�>��u�Y=��'��S�*!�e������ڃ^�����\� ��+��(xuHx��"B�]�t��� ��=7���=�`��}�����1�}N艨�����!�X��<���4�Cd���V���NWz
��=<x�=�6(�p��Z�5J!�y���mą����׈]o�9� >k ��?�t�c�&���7�^�弙"�{�w?���P�)gl���4��`ĖU�;���{�؍�'�5�.ȳ@�}1���a�r��ʜTθ��/��:��U������J�d:CCSS�^A�';��������DH��&��7���[u��5f�B3��a� d7Njw��B�ۗ�Ly��*�a>�p�b�a	J�6����[��cx� 
/�W�fS���͍漂�(��MHҡ>c}���!bp��|d���4�r��s���X�㣦<Ֆ������z.��B��b|�P&/����%Utp,Y�WeNt��'(�T-o����X1����(QYЗ�_ش�5˺S��}�L��%����8����-z�&-ӌ|z8��jEpD�am�zv�-�R�����If��B?��l�V}�voг<o�	��`Ĵ�!C��t��5$�e)׈H��+BH�8G5��{�e������0�A|/'��]���mo��\�� �::���C���ߗ"�Gb�9�k�q�l"U u��5?����=�����+���U����n32eL;�C��d�,Inp,O�����p�JDO&d��Og��gz*����?���A�3���*��
/� ,�k�-�m\��jh������f�1��΁I�,�źh�͸��{b�hU��0-�4;oA�ҍ�8��I�F�����&6�_M���I?Ȣ<�Yi���ڡ8Z��ic�,�{g����Y�m�s>u�E;��c�ЂU19��X�<Ӧ/F���BAf{|lx0��^?%O)�ޭ��#���p<}(�k�L7wfGm��PJô{e��� �<��M��e#�dַ�B"�\����յ5�eK%x��E�+1h��ʺ�=9�u���GOᾯ,=̍�?v^��S,�����;�[/n#ҿ�_��QMy����P�`d��������$��s^��N"�6����p]�ضSh�,)q�	�� }G���P�5r^6�m.S�Hd��q�[k� ݎō���a�:�{��w��e	$<>�_m�]}��OU�P����W�W�Y(�L�	���{z�c�����˲��9FԨ��||�y^k?5�n�^�CCf�c1I���׼m�v8�H�O\����O_�80��L���t=t6;�<��a��AUO��'��{o���3ϔz�Q`=���,:L������M �������	1с[S�̟���ކdJb�|�\�Y�?5��?S��%���=�e��e�
��%�6��X�����~_�v<ŗ��K\�DL$�0�w5M5��L�a߽!��l0���]s� ��8�8�4\�ߞřZ��x�0��UG,  8��q�߳��룅��!`�����)�8��8���f$t�l!�tUڜ1�A��z������~zB�^��Z������m:[�!ٔ:\22�J����~���e�j|�/���z� �w�bg_-���l��b��m��?Q*��ʅh{t��T�a®���[���&����t��: )a�n��)H���2�7ۏ�;��GK��$kR_C'?�	X�I�L��8S�s��u�����A�S>�$��p��~?1Ln��Ӵ�|'�ȋ�	R�*>�����y�t�����{��`��=$̕��VP6�kS��ÿ�%mA��$�2`~��9���q�ػl�����\�>���c����+��A{�iÈ	G�^m
���A;p";3<�f����b��
ت������W�#�'�1Ng^(Ј�x����X��7�/eL�(����?�&S̽��wZ��=�����z��h�䬸W7-%���D�X ��1��8��K��+M��9j�/!��/��|`}�-�j�Y�����4�aB���%B��=3��Č�YzG�:���4e��j �^�`]Wi�h������)
��)��3΀��\�-�̺�	�x7�@I쫭Ρ�뾩��T�]8���F��Z��0��*p�K����R��Ѽ<��qxT��zB_5�����;�?�����᭡Ǻ�g)0,d��WNA��3�!���H��s���{&#Z�NHޞ�uV'7<�\�R�v�
m���Q�C�����#רWlƶ#��K����3��j6��ڭ���+�)�娯�� �B{h�p#F^,t4�<N73"o4������Ѻ�v<g�_�y�D5u���}v!K4^���.�oXޗ��^�߅I����K����P-�x�w���g��qr��m��{�O5F���[.�������t�3z��-/���Pk���w���+�zDqz���%��ԂQ�6�7�G<�P H�����4�'�7�a�,"�GSy���6�ub(ޝ�y`��\)�����M���&�S�N�,{Yύ���(�Sf�	da�+�Y�pnSؗ.ҖK���Ի)5[�Zu��=�tN��3�����6�^w�譭��;��(O4��������_�;��E��)c����%P�ה��Ml�ʹ$녖z`-L۸gp����Ee���04�ms"P���D�Ev���������oI��"7�W�$�𤓂f�?�֩<A�����o�������WT ���#U�0���m��kI�jK�d~DL$�{�ⴝ��ѝ��I�9`h�3��$p��Q*�� ڛ���_�x�N�N5-MQ�]�H�Ɵ���ŐO@�L]�����0��[ѬJh��7U�ņ��͔*ˊo�C�'�W`Β�G`�u~��>k�?]��֑Vb����f�5>�*T�P���Ӽf����ڹ�vPs��#�����a�8�[�t	��{��������֬4�W+�2L9x͕`ʌH^�m��Z4�7}Fr
rvȁ�J�g)1+�DzW��0��A}+�t�=y��z+�J��\��]o
��̞#�j�e�B���D����Wr&tqFt��32��w4�U���{n��n���-b��DOkZ��z{�Hyj �Z�x��M��n&��:���'>}��J�z��;�gus�,�4����� c�<x�L����y�)x�\$0�}�'�g�'w��?���4��7B
^9x
~z�_m�2�_�./Ͱ1��P%պ���K>H���I2���xQ8�^Eh�f�<�xh��&��J�)��Ѝs��d_�����/�uN�>#0�G1�Z������q��)�q�Ҫ�s�e)�'�*��<h�O�.:�J�W��G�;�a��ij�:�CCI�A�}� \���	����>W2,�'4�RR.�P�K�����}����wW�܇,���p�f^�F�<��)T%+�X�h|�)y6ak>^��ޥ�gO,1,	LJ���tVG�G�RQ����^W%Zhe�h64Mf��Q��o�;���Ɣ�^&lNI7Z ���AC��|�Fa����S��:�/{�0��W�
� ~�ϋ�}b�!��s�!P�=��v��[|�`��`$@:5:��>5ʽu�HO4��)J�F*���)���R���^p����ɬy2
#�W*b�xF��y���J�L�����g��ܞ��u�.)H�{���O��A"���k j�7�m�=<!�]�<Áz߯���_��۠���' ������u�
4�C�{Ǝ��8'�B}Av~�X�[��B�<@��Kk������5��T�a�|����x��(r��e䷿J�Gj�i6�	J]�7�D�<�x�jI���Ӧ� ���+���b��LuV��_{�d +�L�i��:w��SA�B+������y}Kh����*R��"�����>E��oݝ��β�Cu�b�kG�4k�T��Tt���(�W���|�&*�藰j��2+�������*�t�/�C+Ӧ0>�2c�:��q��q;���P��hg�|�-p|o���؂�I��QE�A�����մ���K�o�]Xyj.62�ٽ�X� -��8��Wï<cڹ��J;i�
���qy��e����~f���bm������O}OB��~0,�~�%>��_������o]�&B���
�پ��pd��K���5k��<���/zlğ���屺B	h���8i���̯&OP����T�ᛛ���@��Ƥ����w�������+�l����hj�s���I�(�(.������ F߳>a*�I�f�`�8#��YH�u�}d^���T����4|���*���Ӭ�ݟ�]E���?��x,X+d3��,�ְ3����3)�NӜ��g�!���Ř�u�]��3��(C�O��ѦH����:TT*�d�nvZ��-��:\���4]{���+|ց�'�k�
��]ԫg)�1��˼ɼI���b��B�8*�e��z�F�;�6`X��_l!��"��Udg}̽�6���s�A��[~�L�/���m��8l�Q�l)/)q�bX!xG4�#c������*2���XD4�����#+��_M}9G��,>��d׵����l+̴�9��9X4��ٕי
�4��{��F1��i�;��׉?Zq{����.*SĬ�P�V:9�"W9�M}F\�ʛ��Qc'��𷏶�'�0+�嗏���������kjw�N;:��e6���#��>N�J����/�6���q���d���̹��6�7?�g�����d��V,�48��
�@��2�K�"d��_�UU����7+.>^�����\��;Bo�k[R?v��T�����L�h�Uzb�B���:8�k��.Y/>b��?��d��N#��ĞlѨ��dj����IW�y������r �-8�F��uOfs���zm����V,Z��N�r$cҚp���^��"r�k����c�%�[�i;ٴ�������B�p�;�<^I�T6M��Zp��P��s(�߬�;9j��ZG;�����w.�iy���9*V������kk��5�t5���$Ň��9���P�˞�󡞈����S�7a�D�u��o.�]������\��ǳ	��^�;��Zg�9�.rf|#�oU�c:�ux�3�6�3aݹ뫶�J�3+��-̏ɾ��Dʟ���o��nK0$��T�����=%�U4�.��*��Ji�������`!��i�I|�E��A����A�+6O��@{_��(	��O�'�bI<L$���
�hs����c�� ^���䩆�c���6���d��'CfA�2��\z&`a1O�3���s#;6��=o��B������� s��r����"�Y%�X�&�fn���.���شʵw���~���=n�;��>�/��@_a�S_�^���^�mc��c���I��۳����{`R���ς
��S#�ٻN�sv������'邴�1��X��1XlQuq���D"}���sn�_>����3�+�3��9@�;�˚��z<f_W�Jq(�p<��i��z*�s+I+���ň�{�ڬ���Ta�XTh����c"=�ؒ)���3bFF�)}K�ߓ�YZ�۝�[;g�2��k���$�"h���DWj�ʴ%�]i�9+N�D:݀�Ao���W� �F����9m�b2N~�v�0��h�..��Զ& m��{�I�u�8j0�\��=�s���G�r��y�	Q+S���K������`���L�9�Z�`q���u��+E�15r�J��B��0��(B�,�O�M�=��!���	誰鮻���C�ǅ���E����U)�aa��`h[�ʰ����8�ۃ�������B5�ՠ�:[�]?�?���q�`͞���꬞w�H'���+F���C? ���K�zX@�A{?����.��4iU��9s�Q� �����,�#Tɤ3:��٭����<��q?�_�g�af'�����+]�^�
��b�A��7�ڸ���e�j�^����^��醆L�|`��jMPS���;YB`��0��\�~���k��Z���f�M����./�"[U#Y�:晪�?��l{��Q��,���֕hd2�V�����z�d�~�fu�S9����&��R�^F���p5h�0�����)ܒqH$,%0�%*Dc��JK�	�����!�����͆4. �ǜ|��J�7��J^!'B������X�p�ф��Yo�z���b!���MƖ��w�N=���'���yzNU�������4n�����&3�o�O0*�]Ű
0�۝`Hٕ�2̑>WF�~no��z������8m�D�-cxo�d����>졕<�'k-�p�Q��P�;�T�%�5=��j�a�f!@z�����s��ρ�j���s�peNI��k����S"[���u��1lF6�����UQo�5�*'@�I�۱e�M�8	��Gf��>)-���s�/l/�}��+�i[�A��m���{ْ�j ��?0�(^�6�Փ�+��fƞA�\$����@�)cU����"���Ƚ1�׏���A�Y��M��{{��w��&��D=5�n��#��mG:��=Oٙ�A��J8{X�"�X��[�o=��e`��:��]r/���8"w7��4��QS,��糟Vt��]�_ߞ�����hD�S������1Z�D1j~���ܭ}v��=.��Jw��=.�T,�#��J�����F>`*\��]��u��-K�KB��y�m8��Ҥ�a�A�µ�͋�E���;��0V�Y�Ã�R>�������Q�K��a8�,`0��  �9g�;r��qW�H08��\��㹛=H,�+���������(��^��I��_��߸Z:p7�W�ú�����-��q����1�1^�*�I��7z_a�2��*:n@����H,��9�s�{#�F�[+�����9������ػ�UuA�t?�$8#��X�DM
�	zG�ɽ�=�#.o�O�;�T�m���'C;�vO!X���J[��H���E[�6�bf���|I�	2��3?ECz�M���.�ϩ_JH�%]e�R%�e��Ba��`�$�r�$P�~[b���>oO=�����F'�Ԕm��㠮T�+!iAb0gՀ��ӈu�;�]����"EL ��-f��#��$��Z�ݬM/mR_�(`-�2��N�zC��}�R`����،+�G���qeWlK��Ub:�B͎�Pi;I�mT�F��ۚpZ=	A�@c��q�WQf�җ^�?����4m���v�<���k?��x�iԸ�-����/�H���y<��D{���	��t@�U��6���e[�����\�hj��h�p��8�Rj�W�O���iXTr�/(��]_'tp�
+wm���ψNZ\���9pU���u�l��c�H^�餡��R2��=�s����mK�m��X�+��m���疸eӢ�7:��f4�%Uq�r�����sF�zR��h
A)���
F����-"�A���+@^�����GQ���q��2�Ej{�E���4qE̙_�F�{n�z.�:a��u��c;�mH���Ժ��K����RG�@Q����2����5���k��iY�>�
��d��. X�P�R߱z.����L�b�bZW ��~Z��h�����?7�d�ǣW���y`n�̿�w��`����N]#U�b�倥u|�Y�*]gD�ҥ�xh�z~d�K X������i�|a���Dzs=^�j�>Jv#�?�b�5"͎�0�*~X帵/J��e���2:��B��o�(��۠#,���H��q���7�W��IT~tç}zV��35)�?Mk���F��'�e�I�B0���ށ���7���J��Zh�h{:6�2<=�����g-N3�\������'I>�	��1���'
����)�~����~9E���Fd�guU��q HL�Iy��3[�5��"����E����UN��8羛dOh5��`c%Z�����e"k���kt�)�YF�dֳ��7ߠkf��t3Z�l~JĆ���7�x������/t5+�L�#�L5*���(�;v|��L�����'�d2���3���l2���+D��{O�"�m�RAg��wz��wD�u1M|����́;j_L��:�jeG�VX�5>+�Κ���ez
l�Q?�l���˻���DO�͚f��
}�&&�6��}���E7#�3�d�`薗��㴖e�n~V�� V�R�ʙq��-U�����o@��k�"���[iTҚm�ʥC�QF@�'YTdeU!J���>w��E�����A}������+Th��uN%F5�,Kn_2�]���t`� U�!��瀆��-�	�(���,[�i��p�!��q�*��O�̒o5\^wQʢ��Ɏ�\���N�]5��U�,&�zB�R���र�H��p��R;L�����������6°9���~��`����Tj*�.?^Y��O�}d�Ӑ24�`k)�������C��r���8q�;�Tl��U�X�G��5��� �	~ t���\YF��8Ȼ��w=n��#+VNRs;�:�} +�ןuQ��J��F�X�ľ���[�o��j�K�|�4��5�2��{v����4؎�ߒ�rW.�U����hw��z�mlޘ��tM�F��[P�/ʰw���'���G��,b?��X�7�/M ,)��a$�%�b����d*jɱ����1�����&��H�J��Q�)�I����_��1�����;����>�zQ� �y���hT4�V����'���(0�&��з]�P�s��㲇�0{��A�T�|�*�Y��p��.d߲�@oF�0[	���-�up-�hg���_l�-�k�����dm��h�(�?��;͸,{�v�o#��;�xyw ����l����-ם��Q̝O��n����Z�Qb��TBv �v8;2�A	�/�M�%_�D��:�@m�)7˱a�^+]@���K��`l�v�"淏�iC�}�f�R���#B�ެ�Ւ�e���}�^/�Z�l����Qt�H��]1����}S��b4��e!,.�[��vl����f�h���h�y8S��M�����|[-�쬻���[�h����r�w���a���g�%Z=2�C�j�سI?&iZq��S���4��*O1��=��L+;-��0�l�di�t�thEo�K�g�6�y�ѰC�=>���؄6����{�h*E`��RU����Q��s9x������.{:���xNNXB�1%<�#�P�2^�#nu��W�1�6-ln��D�4۳ɜ�_�����s�7&���	�?���+���C��֑��p�o)t��{����("��s?�O�K٭����4���-:�.qگ�[:8��؟�4S��Γw���f�p3s�#	�X�[ d��a;�	݄$dA)��w?(�tI��������%kq�]cF-���aIG?��Աy_956.��E����ed ���K����ٕk���
Jy��!kǚo�-�vZH̜蹊�F�fr�������I4�k�� *�2J�6�;e]ɠ���i�4�E���h�m#���Ț����t�����x~i�p�a^q%	�������d]wn�+Xz��5��u��}�'Y����Q+��QL�f�(���(_q��NH�L�H��BΆV�@6�HQ�����h,h�:Ҳ�0(�8�*:�:�KH�=����H��푦Рw����I�-�X�*��G'����H�����M�8Y���f_����B�)�����ܰ�3Ӿ���"��5�ϫ���/��J��oqc�]�1SM!����s��Qh���mY}��}o���c��`��͖�%7�}�V�u��������C~�l�����.=�Y�2�99s{��B�Ci���xE�����$3�dg]F��V��tG4�K� }��$�q\蔰�?9hfU�~��ܾǛ�A�4�5�x������=�\���*0O��0(��ٴEzgׯ���	���dj#*���1����pi�|Y���x���md�zh�ϿHXP~�8�פN��G�Q�C0�A�=�G}�R�y�8�q����A��T6,ds ��OCs��ٓ���"�8o�yo�>������٠mk�B���B	y)�p|VB�����?>�(�� �M�z��2�VѬ��V�O������[����������ewԘ�4;�W��}!�V���Z�|���� E��A���	ڕ�	��[0\���{�W�2�<�-�0�?Ӿ�,�̲�w6lv�NA��@/k��\����/kTE�5
47��=o[�=�[�ݐ:���<*�mH���DC�L�h�2�sE�(�s�70U��*��,�;���/Z��gu���05{�2P-�S�D~8�%�N�
׍�j�F`O�cJ�Y���9w�e��7�Ԉ�绗\�;0��ݑ#�+�=4yd�����n�,T��@��yM�SN��F�F�od��_d��ob�pפVs|�������]qJ�O.<&�Ԫ1�N����VV��6o5u����k�m�b*u���ğt�	����KC�A/l��A�%�w��.��܊9���I���~���lc���w4q?�h�IA"�	{�E<��Ѱi�)`�>'=aEp#�0�gA�zL��g����F�܄|����]y�O_�Z�J˿��r�8mY;�M%���o�y�M{.1��6[�h&����M����'�#nﱹ#�*Nm
���\��	7�_Xo�n��!iKi��0��;��Ӵ�a:�$|^���z� |�Ϸ�U-^xM�i��H��z����")��4�X�����g�-�wJ�M�W^jK� ��zȓ:�ޭ9-���Ga�����G��4�Y��&M�e�7���ؕ�e{�����w7����5���^�3PvZ	dX���p�O�φ
�����n��8�l�[�r�Ժ|4��ފ1c-l�=²̨߁[���,ñj¾j�~ǝz6Pd��8ܸO+x����	�g�8ri9��q���{�����6W�qM��I�:��|ָ?����<�c�ǀ�p�y�^�����m��u�k������_&l3l6t=��<wwX��94�v� ��@-k������Ѩa[��:B�\�U`�	��jrO�C�ϦƦj��wMTw ('������-fx����lǑ����:F�K�=��q�/|~���{����4b���E}�U��&\��%c�T�BT.Do�\�cvUo�7�/��QwT�1��JL����gu�G��m(���J"���5���c������F�g6�\5d<	�s�#�|~]��5���f7�Z�:Z���7�2��jͶ�x�-�D���O�w΁��o����{� �E2��H>�|$?^:=y>�:r]-�ހ ?��w2�}-�*��U���;^��H�J?:��9�z��p�t�s���L��Z����E�mf&�o��&�ǂ4T����cJ��V��(-h?��W�4�V&���;�OM�����_��[�i��lq�<��JD5�`s����qD�Y���fɈU�����Hͻ�#�9��eVT}<H�$@��dZ���N��z�������Q�nķ�v��{cHQ�TV(��q��WB �0��.��Ǣ��*w�A�*L$==�Y��J	σ�F��/A����*�8���o;^R��^D�n2�̇�_���N��v,�]�%��+a�4l���E���{�P
"㑣���YeC�ɳQ��'t(��f���@=� ��(��ѵ�P}���}�Q�)K�O�q�x�b�~<����&����B��������Ɇ� ��x�`�D�_��c�^�i��n�G�F��LF��L[~ǁ�����;r8��j?�!S-�\���%"�u;h���_~B&S��M�p���Xc�d�n,��V%��g���9z&8.��Ϲ�t#<K�ɸ�+�u&M�����3�[����G�8������l�F���t����o�-�otv�<rs~��"b��JpS��/��Tt$]�.�1����]h�i�|�M�5�+"ݠ�#�x��q�VK[j)t�5�w�Uwڨ�!�K����#�������]�zk��	�N�1�g�7:|c���׽��I^����l�'�WS�ʔ���N�ӄ)�����n�5ȿ�*�����p��z��+
�L����닎;jh*䰱�e\g�)�Ύ\��_D�	��d�]m-:��ԭ{C�,$����;WR��^P�)�HQ���1w:����O�Ō�Ŀ������7%��P�x'������������i�[�c����5X���Y3@9^����K�Esß����Y�#l�L#Ҕ?�6��s[䥬�zG���߬�E��R@оqΔQ9*[{v����1Ū<�;�S_��|ϗ�0���H����E�	4�Y�N!�>�}��o�ɼ8"킰]��w珏a�����j���p)�Hiqwww/�Z
w��EKp�xq���ww������8kVdd�w��L2��́��q�0.�0G��n��<��.-��/����[��[
�;3�c��\:Z���V8�SKN8�z�O��E핲�gY[�����s��QBI�in@���1�����%�1���3�"�����ũ*�]e�o�>	�i�ՠGk�����ͺU"z!�F��f�s��T�j ��F�PW)�����G�K"JSl��3�����
oB-���ٓB�5�:���$Ye1k>Q�@�I���^x֓�0�̓ܶ{��k.n3�)�2x�㥽��=�E����ʛ"��=\/f5�:3u��B9�������`���S�j�E-`ϟ+<e�����P*���j�U9����2��MP�s��W����!
r��E'��LW6]�Z<�-^5.A؛��`�Rx�f]��l�L R����J6 ~"�WIJ�ь�)[��1�j�����e��p���>MW���K�����&J�ǌ��ƆXK��ۅ)+���+󨔈r�~���n`�8+J*����lcːi��)dS��(�� =f���9�E��Q�ްDd~�2E��B��$?�/�x1a���<�# $TH�"�4v�f9}|��e�;����_�9�>*��FzC����"?����%��x�Ș�w�A�<B���{�c ��o�~-�#�C�5��1��x�~=o	����E�'�tο��M�Ï?��*�L�@�"�7���s��8%Ī�Evȸ~�_��G�RG���S
���*i�׳ȩ�T�jb|�s'�sP��	��Rt������[��V<b�-��(������'�~�	P��$3��p�)�m+�օ�!�δa�������AL=�nm�a����%+��HD�����G>�_zj�.����l�ۧ���-kD�NqTc$��Q�${F���S��D��ҡ�
�t/�6��rt6�}O�eǢc:�r�I�Wˑ�]�83�{��l�,�Q�Z���N	s\!�-���I��Ĭ������4�Cx �-���ǹIG~�F�*�7��W@` T�j�m�����\w�T�qg"E��q�+!����
�t�s�2ׅ��WBR*���â�"���S�'U��B{U�p��#��!����'X�M�/��T͒E�\��c(�:ܭd�*eW	�fr֩����B>m?���/�0����s9$a,�g��,�m[����_d�㉩zZ~��t[�ugE� Eib���_�������ʅ����T��M�RhD����ۢ�Q��Ǧ~�{�]_D.E�}']HS�f)d�5ִ� |Ddf������Hmy����J���֚'������H(/���V���d~^^���Mϒ��R=��nq��D4=6E���S��/5X4��-�8���A>k͎��T���G� ނ�bE@���]:mƓ`ޭN�o�)E�o�,k�V��hg?��r�Z�A�BM+n��Q���P��0���ت�W6 *�&{۴m�닆�BU�����*�!׻�τ�Z���V�5y_��7"q,yｺ��Cr�%ku��9�r^�v7�!����t���/�%q,�rq>��4�_{�f�4�LGrR�R��a�zK�^�\R�Hzz��H4VV$jĝ�)u��1ʼ��6�H���9:ed�g���u��4������JD������åᶦ��s,�2���J��������|��Q��2�R�R��ȑ�u�AS>��
�C�X-�SJ
���ٰ��|�������-cS8���bC���Wׯ�ٳ]�^� ���~���/��|��j���b��yhv�W��^�����Q�y�+�'}�3�*c�q�q rv$q`�p�7�F�O"h�¼����r���G�QyxT�N��p�?��\mI�.f���e��4�g�*Q3���9�t�(�}K,�����9Z/�(1yx��P-�xF;o�na�iN�b6GJ����.�	k+�϶0eĐ[f��`��C��|Dr׼<o�\�"0q���*+���0����7�N���	��U���!Y�'�j��'z��#C�����1�Ԣ���ޖX��tN����?(n�y\�-n��8q��
�-���!��zP�C�\!�����}g�ԑ�Y\4V���pa���F����@}B�Q��4
mB'���4����:���&�/���?��iW�w��J�[������]p-�&O��<k�����穗�D�>X�����8�~}=}֮'^L?��rqC��t���.8� 1F
���P�y���;�{���y�n�;���qc���g��k~~�`�����hT������m�D���M;YH����+����[J�/w�A�����΢������
���.w�1��mL�?�5�c�=���4b11�)"C�&�Y���}�Zo�Ľ~�Ck�ֽ�c�mq������ۘ�5���Q��4�	��w�m�.�� gZ���t�I�-��u,6�d�טּ��5�?U�$*��-$�&����K�bj�G���v3��<-K����L�>�c�m\�n�,�R���A����\l��cJ#�k�OOM�CO�"�B�=yW��K|Wڒ"%�L���[�>l�-E����ɳ�#J&�P/����o�/׵df#N[*.){�i*���z���Z���d�#��n!��1�,+�u�˔[�#N���}��7�aO�=X���H}�	a�E�	��}�'ݐ�N}�󔍔�)�����^[�����#nn����D��u�v S��w�v)��Y��F��p���~F�!8I�(�j�������hJIb��FG�;�ĝz�_�,V��n��NNl��Ϩ_P��i��X�їyʦ/���Z�;.@-t�G�6�XN
�M�PV�����Ds(K�6GR�#��#���^�lP]���+��G''�{7w����܄���c��q)��ɸ����$���+�A=ޟ��\��JſgNuc�^��aO���o��KÉ������uՈ���˺-�ΖdN�n�� u��Gnd��c��[��p�@��� ���p�K��e���
ja�G��Wd�u�y�&���ph&�gk{��3Z��?P���sEֵ�&[Z�����e7��i�����I�AG�����E�cf�9�^��د�'��yT��l� Ժp������g�H�z���)�;�+l}�;r� �LT�<B��`����_���>��Gǧ����~����641��>��><�Oؚ����XW��GK�]b���u�Hby��e=�9E��y�єg�}�ck��B�4� tn��R�˧`��4�����IA޶�:��8J�s؝Ne��\�	�zeKU��z�P����Le.�1�c��B��!�$��=	5*�7��nI���B�0�w
h�@?~�2w�!��p ���Ƴ[�0����fUU��`�Q|K���ްn��#��6mtfvv�;��fS��kNa�����J�E�`�<����ǂ��氠�ɹ3> ���?E>i�������:��n��b�ѱ=�D�������^gr�;>�_fL8g����2��]W����R�?t��6�N�!
E=�uV��S����I�ٕ\m��N����4$��'3���g����v�������..�'���ִ��ԑ��X��%E��&�ZJTʖ}e����z5�L�HYo�H84����Uz�y��GyJ�ma���q��]c����~�q�)�]����aF���Qρd~88&P��0��_�C���A�ڰ�MR��ȱ��O}��՚���� ��=�������nn�� ���۳��*JhB�DΟ��֠��%���+�}	]V.?Rٌ&^��Ox]��s�P�t�E���7���I�~+1(�05�����5w'��� ��j�t�%6�
E����.����?>��i2��5�h9�$�,��%�f|�F���N^���J�����=��]��'PIkyTǋ!,-��ϋ+��q���֙7�R������\��(��t*bj��M7�0$pL�86��;�R��4ƮF)G�����x7v�>$
4���C;� W�[��	��n
��&��BV?��� ������ ��R��U���OɤUa>)��`���>,Y�����B����F 4u ���є
�4�/�2�%@	{����&��%�}_ <���y�ѵ�z���_�@��^��D�ad×M��ܼ?'yE�6�����,�F��Z=����,�_�l��E��ŀ��lP��c�Yƛ*���J��W��{4�O��zs�}��"zZ�������������:��=&L_yaτ�^
���J������-��#���H�������Y��sk��y�D�W�!y���2S"E�@j_���z����`�Z��R������e��0��A��-�nY)U�U�7s�ZX]"�2�YS�5�.^��a���&�-� �U_�hw;��b}�ǫ��\��c^�9!Y�f�)�fgbsj^�����h���P?����r�J���
����sC��@�9.9��6��Ya_~ّ�.����ú
°�h������z�G7�Z�-��2��ɗe����/伨�3�>����7���jA������mÝ�k�L
:���{L;~�`u�O!������AΫ�̩��xr��:jd�>'�\����`I�t?ҫ�]�6�>� �uZQ�M+�3f��=�"pӪ���'?}�1Myt���e	Ahj����#�t���p�~���m0�g��D)����С�rdM+)(1��&%tT�2��0\�E��_�n�o��t��p�O�L�XY�,�`ȿx�P����nwc+���z�&����pA��H��kd�s�+O'ķs��*o�����
�5'���������B��"�7����?d1k9c3R�9��ffl�˯���A�����-Z�u�7��)�$�ϐӾ�齆᯻]�@f�vf}j|�����G�|�ڜ������V�X��=�X�ԓ-P�+{f���'{="�>x��|�|b�x�c��|��{5�{>x��}:ʽ �>wT�<V�~���bv�?IXUR(�j�J��DeD��a/��֨��Y�豔�7��w��U��͔Kma�:n���9�1�%��O[Y�i��Ή��Qu�-�AK��z��K=���6��fL���(�b�T7��:�x~oE�qp7�+�)�-�����T������g��>����K����LI�~��}Ŗ/�^#M�Y������!'#�D!)I���7Nzwagt���qFl8Hj���=yDz����S˴J�׆{��� 25G���}g�k���P�?nww��l:ۖO��f�"�s�-$*Y;���W�a�D�����e5��W0�/�I���Lwee��ӔHϠ�ܾ
��c�Q$�,~�Ƥ�k�Z����GW���m��<����: ���^���Q��1"'��uύ���6�D+���mC�0��xC�[��*6h�쉷�f�%|����@����5�4��#��+�*��8z'v!]:�aB��w�m��ܷ�5S��?��%���}Tx�s9���"N�E'�y��U�2e���n���*;HZ%ȩx*��{��н�6@Po�^.�d=o˭%-
WY�V�6$�CH7/IdI��<�����"(���ފ3*j��z`��~I
#ck��V��)ID����:+4&�*��I�{RZ�Q'������8%ZI��"���=��� �a���+o��д��x�W�y���u5B�H��ƭ�fVF�BG����h�=o��pK�g��aҩ���7hn~��+���(3s��Ż�\���/:�/�ܗ��9'mtZ�x��&aY5����k~}�k��b�"���>�-i�8#LJJҴ�����OD��vM,��#�����=Z���s�������O߲���d��#g67(a�$g+B��8��u^9lrR�G��|�.������4�c��^IwD
��rq�P�劾8�x�/�<-�+-���ܒ�3�\?W�Y2F��ޝy����T'�Tj0V/�[�)�DP;������7���ʢ"��Z^���}�ós��	c*�T I"Ƃ�-�\S4^�:g��2C�*��R��ado��~����io�#A��%q��RXu$۴Ŋo
q䢠!R���݁#͝�ľ Xa��XAud��|���a��)��eC3|�_G��@1"^���jՊf*Y~�S�$,���E �����iq��^�H�֗���Ru�{��?�� �iG�P��m2,�


�[���Cagg.4��#*�w˷��)K�3G�(�]�&[!I�D������8m�]����XM�1���
����$c��J�@'1X-ݍu�q��z]��w��NW{c�V��|�������ĂC���ҁ������hT�5�z������k�3b!�mv~SSK&�� �ޏ:�����߫��$�E1�pQg�pM-��>Yv_d��&�DFz�,_��+@�9{��]���T=���z�QJ�.|��5�f-��ĳ����9&nn���?������o���]��A|�\]�/��0��37�QV�6�j]��Ӡ��A�>E�2�����r��?���C�--��}ggglb�M'=�"�ܫ�܇|b+ v�D��h�냓O�7����٨�\�R�.A���%��i�����j9�����Qo~���IS�Pߔ�OH�_]gO�;7���j�����)&��(����U�	�_c����>{@A�L:� �����"[�KB����ﻵi�BFU�#�	�I<�t�9yxz��:{WaW��AzVF�2*����5Vz��U�
.�T0���4��J-�cLO_�������N���rk�,�w� �+B��="��V��L��⮇��jA���r��kQ
珜�oA#u���X���\���ߐ�����n��G�wĳ�x�Ҋ> T/�T�#}!d���g��Px��/�s�&���/u�#������Ul�
�lk�;D� ����Â�vx�Z�Ti�-�MQ!��Y,�'��W�
��a��LQ�2�ELi^{{���h]��ں2�ڇ���c,��$lÊR5	m��"e+�������A�)|���.�p�`��W�3Di�t���a�K��,O�-�*�o��u���&�y����PlS�9�r�0׾fA�],��6fQ���8(l�5p�t��fy	���,5�X��	7H�[��*�r���ˍH[h���' ��^!�j6�I#R��_��ߡg�������c�|p��r=!�1�s��m#7s�"��FM���04K�3�d���a�b�U3�T�63O���z B�%�����1�l,q�Ff?��;
b-���
�R�"\��m�!�r�3����N")%���s�������
Kz[7	?�ة�/���'�b���
ڡ*�f�Saԙ3����;��FV����������n��_NA�fqĻ\�"��h�]�BYk3K�P�7xG"��28mvE1X��-��Ӫ�aX("M�"o�l�5�U�rV�Z�d�0��j���-�2�gF ���V�K|�~�}���=:<5��HULc�⣋^�6J���bK��em�kRt�w}��z?�hrd�k���f����f� [�t�)6v�Y�މ�%����Ҷ�������c�!U�6�۽7�)�*w�;���> 1|v�%�=Y� ��9����
�U��F� mbFc|�?���E�[�E�_�!yF姂��(13�b�[���.X�n�����k�5�7͚-Q�<��]�z�����6����%��gu�i;��`�6�$�����X�Z�kZ������ٴ��S ���p��+E�	;�v$O_>�����0����gF��:`�����h��&�IC`k�?��/g�Rw;zPfG�a��.�]���E칑{#$DU�����$�����&s��؅�Fa
�vDܵ�+,
��(>�|�����`��G'}e,ɉ�cFz��a�Q8ӯ�E���15�6@`�ʑ���;;;�W����w�箫��K���as���]��I�!�h[�_Z��\�"�{��V�x���F��Rc���%���3�/\PP��E{9���yչ�R-<�	��:��C�9^s]���8�z�DWs+�H�ɗ���Y��*��>�iH����UY�����Y8WIPy�	7
��ƛ0!|C��'��v|b���(/[�=%[����K&W��)����7w7�*Ec�f��y�@��E=d�f�Rw����,,�~�Ĳ���{ؓ�MK��kȹ��x�?~l1[�]�Ѓ�]@|��;w�^���z�'�T�'�j�z���.�[Y�+��qa��B���'D�R%��k�{�r;�����	(�Η{'�~t��<?��^l7���#t*�JԝL+�m�/�ߗ)���V���N��5گ�t��6ú����I)��N�*�wIx��xQ��`:Ec��2E�ٛC<�7�H�_aњY��7��*)�R< � ��#hmm���޵K
�M�k��bd��;�r��T�Y���� *�^U�����l���u%)������"���$��_�֖��-~�p��u��RTZ.2{9Е��u��W�T�d?�؛yOZ'c~�pN�`��	���șW�j����_�V��m�NЧ���5F�"T29�+@*'ҽH�d�B�=#�]�ho�T��i�����l�����_��t'ѩkmv>~Y{[):5��&HW�=ۜ���"��P��#!�٤U�����7��z�
)8���v��\:0Pl���M��O�+�glT�E�U��r_�a����:���c2J�+!�� <�s��^�<�nV�
c_n�;�.�+�]/��R��	�MZ���"2iW��,-u��-VҤ��!%���=�����7S��'�o�d��b��A,������ӭ���J�vd��f�7���~�:���<�UU�e�����'x�[�k�z����?L��{9Hv���������-:�Ù��璞�G��2�H��� ���m}fb�+hW���6�X������: ��tb�9�69��6����PG^�5��9ƔB�]f������@sW� U_Y�Q���_�8�G�܀+��G��>��ws��|�"������~bfm)�z�h��w��(H8�0�w�~��w�,=MoRg��T,T��]��ĉJp�_�my>lxv��]��p��t�&�i��		�WR�d�KaZ��;�.����*o�ļ�Ia�qrz+��JT��/�4��ɳU���bt�0L�YF��2�F�d��v�C���FSYvo�N�!1uq�X��(��*m��Pſf��y>��Q��GK{� #k�yb��ECߘ2��Z�KY̧y�$�.59���d�����@�A/wM�g��?A���{<V�ݞ��>���������EY{NQΑy;�y[��_0����?c��㭉J�`? ��llR�	��6���nNj=��D;~1D_2��s�561���E�'M���ާ@���������!��1�����,��B��J�(��m�Zt(����`�d�����P�gа��d]����o߻.J�LQ���eE9�����%�^�=E���ݪ���D(G��*��=*��;J�0��[�x&�N�v7I���y��� �il�z��Z'����^��}�s����0����;�t�d�Ί���e���HJK�b2��e{5��v4�wqb/��uO2X�,�nq��Ly@*�k���[�rXm�|!�D�{��VH�˼�Bf��lȻjq��
g`�6��j�j!�I�n�<=����N���j��h�_�j�L�f3�x�3�,ҕZ��֎=Sdl�Le����w~�4#���� %zk��N������4�����=#R�5�&�vf%eÉ���^��{���Y����(�6+���L�a�V�Z���cJ��ʘ���1O�Qk�+���1�^�3f�֚�����M(i�~,��*t������0%`�b6ۻګ�oI�[�������u�SW�0"OR�
W���\�`�I�<��S��a�����@zg��0^L@Lh��_���]�H����1S�Ո��,o�	�#�x�ɍ<b����a����-"���u�5�Z���T�ݾ�����X��i��Q�����{�5�4>��ep�,���tNqgu��"��-a>��H��ۡ[m/�*9��CC���ް�4[7�%暣m����7��I?I%'_	���'}_֧]Β���kZ[
q��9�Na,�-��]X��$��0������&t�%�0�_{0�H�j�Im�U�~٤�x�o�|MF�j>|��r.��II4�.������V���j�4`�5�l�j�o�+w��$g�zN�6������\o��]]�h���2`� |%��a
n�g����tRe�eC�>��F<i�f|~guZ�/�*��/] I��#��|����Na����nY�Xoݤ�����܃���7��X��>�*�;��4��S�ā(D@�rXVi	�]�<�ӌ¦�9`�iy�><tv�=��ݬ�N�[nи_��y�M�nvf�f�cA���j�n-էM��0�<=��~�OLL���3�ߦ/Ա/(/�݅�'���UèRt��=S�ϼ�B��"PM
�qWW�D���ӓ��5{��9�hτG<�x}y>]m���� ���w竃/0��t+׮.�a��u�� �	{h�ѕ�bZhsGg����cX�����"/׮,���i�x�����l9V>>5�Ա	K����xl����u���A�(GGG&0B���D�"�w�:����ߴ1��ƋQ���Ԝ�i�+��Yq��E�����F#���kW��9��=<�O96��Ȍ�����F�}R٫4.�+���7	��tI���g�z����T1��iLtA�_�,�+��FqpssS������Q斛^�*��m�~��a�u�ׯdxlF�`�����~;vF{چ�~�������s��m�I2gh5�2�s�n�D|�}���������j�Ny �{�#�hO��U2�.  �e\7�Y��'�����2gzt�'}=�RM �'ȕ�MzWA�I01(o���4m���=��u\���V9�������ш8�H$�܌6k�J�I34���bq��;� ~��l��_G?�yt�������z��.(X��#.u�� e�8˜!�6`1�a�c�)�*��h�<ߩK����R��y��>B�e�'oK�ee0�{� �yޛ�[NQމ�Oi�.�����{��u�#g30��C#��J��L�a��[\���#׌��t+�����ﻺܽ�\�TXٝ]���f49��K�y���U��c\EhF]F#���2l
�伹�Z�F�Q�~������a��1�'��'���N�;q٫m�\�u��5�3%R4�ⴘE�BWVÇ�Y�o��H���o'�݋���%8�j����J�p7,��ጻ!4����-nG(0�`�踱�#�K������Z��q��Sqc��R��Z�rKk�p��0�qy���<E&����x}����e�9��\�e��6p������������d��𝖎�A(���������3��������r�	�8��y+�j�5�7�y9����u�쩛�1���(��t�D-�@Z3C���K;y��;�
������ַpXmt����7w5u>;�\��¿^�^��/>�B���	f�`�U �qG6�]����%�{Q.�ݙ�D���5�u�Y�=��=��^�>숽���^�_{_!�Wė8�'ɗ���ɶ�}=��,T����=�iDI'�j%���&����bf5��1fQx��٧��(��o��r�^{��yOo��^��Ӿ�m�^g?�e|���������_���J�3K�a"5E����qC�2��s�!�m���@��|e�
��/��JN�uon͛	�%��w���A�K��):g�VLE��9��lui���L+`
q��� �4�ml|\�i����k�.��|��;x�B�:W%%U��O-��J��#I<��?ş��T� ��@8gL���˞�2SXg�A��HkU.1���9�oI߸{�bo�*B'�8#�cف^h.5��*���=��;p��P��så���ekQ3�OȬ�X�
X2�"\��7T�'χaՀ��%~׺:%e�+X\]<�I�����`oT�sIL�L3ѽ1�ouy^��Wh�6�d��KTT�H#ϰ��(������i-�O>Fܦ���Zu��:���B/l$�:�$%%CՇ ;t^��x��b����c�f�ckkă��{��gV���E�sf�o���t����XK�0z<����#��HYDk�({fT�2���P����wq���2�|�
��L�������G��qV��w�Y�p6{5R�7�kG�.ɇޕ=
V(DB���xz�4${����8gg4Z���o�Փzwf~i?m6Cd�Y�!%+��.nn���hiA��ߺ{�f�����`%���  2--ퟬ,c{���K����"A��e���}˃RM�w�u�(E�a����bTbh�SE��O*!4��RI��ϙ�����:/�o��e��=䬲��v���#cz"|
Xy�'�m����2-¯����h)��'/������M_�t�pM��){��\��n~�)/ �����iOp�__J.u��CE�9k����j�y�JQ%��}���qǬ���_��D��E8����R<!�?�,##�#��m~<6}cG�T�v��;�j��oV��P�T}^YOO���vl�0"l��l0��+��0[��Q�5�m��p`�+)>�ϕ�R���߬T�:��9��fuˈ�X:'�|E-G�3��MI%���\DO�m�H
&���!:�	���:��	���혀6;��Uz�zz����,Q�ȤU�S�O{D�5ð䲚�ك��=�����g	�G��w��la�V��ZB���gWfV��T���;�(Q�\J6�� �^�F�����>��\�ztx�#f��e��tEP����3��,�#o�Z<)O����������J�����k�����k?H+hƝ���}���Ŏ	�Π�Y`X�����+cR�&����2+ӭ�:q��ɤ���2w���T���]m3�\
�z����j��N9�|���'?���{a(��^���z:��ٴ��F���\�R� �m��ˊ�sg�Ǆ����*��Y���c鶸��f���3Ҍ�x��oM]�x�{Ĵ�$����	\��6��ʇ�b�2�ۡ�(�A%��MN�mK�d���3i�gf����ep���|.�� �6ՍQ�"���<Ӟ���?s����nllljA�����t	�C�WkoM&���F1.�ef*�B�j#�"�X-�&�_W���I{fyp�4��zw��հ�o�)�`�Qw���+�m��[����#�q��U2e���d�����~Lŏ�X}��W+�-ʴ	#ʽ���ÿ�������0Z;�������`�
�ʢ'Ú��-�>��}QLn	#�A\�;@'�7�ߢ�v��S��q��F���YW��K�[O��;�.8��yz=OQ��[�����>I�VA�^��^"�^fŶ�^��/��v��]υ�K�a�2~xt�W9~U�0����70��^��<;�E,����L������0�tz�l�}��t
H9ȁ�^��
CR�/�z�cc򦔔�����AV?�b�/*h'A fAs�ZS�Jրi�"ڏG��p����?U��S��c��,Ӯ��t�vi.#�,g���'^�}��ϫ*�6x/lԴ�9�T�����IO8����� ��Y�3���b�/6�4W��� ��oCM�i��_���c��1���:dZ�g?542��#�!2s�}��L���qF���U�^�84��͢�x��k���4�=�ޮ��l��y7�K�j|�����ƕ7���U-h#f���f���0T!��w?Y�^2�����z=�5yQF':�?�.8�g��2���j�y��{=(T�ٿ��"�ໜ����T뿯_7
���5u=�p��KS����ǖ4��H�'����[�/�0���P�c�Ml(��!����袈�Y�
�M븡	 C�@٠�(�'��o�LM��DJ���Y��F3{�|�\��}E>9U�"8a�Am���s��Z�8��|޶���j�,���CsO�{�mp��]\�;����]�0U_&����>b�=N�y���j:���v�v��^��x����Y�(G��//p��G������Ɠkw��>��z�ņv0\O�;��8�iz�����X@0֠��U_YX��o�R-[kl*�� �Ҫ1y�����+:�^��]X�e~ R�3�S����i��:D���lbv�-0
l�,������K�D�eM\ۓ-��ݘxX�Ĝ�kk&M�T��XRR��(����]�[�����_�����;C�V6oJ�h��k�����C��0[<u57�q;��!v>�I�,�[*�j���w���o�&a%΀u4�+:B=N$Ģu�I�\�-���f)H�T��Kdr��;Xџ��쨬�9�9}�0Y������)\��P�&�f�Kܗ��x[T��<��:�bX�����|���b�þl�ffgG�</a{݇��?-Kf�_a����pwߑ�g����SZ��Aܪ>�b����_��%�q�HF%�^�n�M+�����sXL�� r������+��.*$7Owdөs�fHW;1��_�P�O鰖XM\�'h�k���*N��et%ôR�/�-���'S��P4�9�ó�)W8����a)���"{���F^�4�0��,�����w�&N3���$n�C�6�������̶�c���ꟇSzĂn��B}���y|�%b���P��,���1f�P
�/Ӌ���r-*�i�A��X��8��j�w|�l�&��SZ�SVzJ�3�ԣ����~^��l@I,����R��;_�%>��/�f���]�`���K�0��{ �Rfp����d��.��Q���' ؙ�c�,w_Y��Ϫ� �	�����6��A��J�l����H9A
�NQ��:)�ܷU�$��&ʸ�P(
?xHV��'�;|pU8Ð/�����i��9�ۙ9���_�S|�>4:6�C�W�}�c�i��V��dK{�=o�Aѥ~��YQ(�'�m�䪅W} ZBM�GՎZ|���C�܀���{�C��-'j�7�V�����u����U�ĂA'��Y��R��#�&<(E�:�!��ݵ�m���ۍUv̒��!���"o{8��'��������	����Q��[�^�c��G��@DYgӗt\&d9����Қ��W�T�y�,G�#��X"��$�����iS(�&g�.��O��,���nl~�����s�g��ǯ��P�|�q���,��Ox�켼*�}�S��mט&,2 ~J:��o ��[� D�5	�bmy_� ��c~7}q��z�8�M��$:,?ֹ�1��%Vl�^����Z[���$�Җ-͸-H�Hq�c����)P�[�|�=y[5?:�V����d6� �A界 jɥ��\.�ΐ%����T}��|�š/��dq�]������c��X�ʴ��p�!P~����WC�O��C7=�����h �3E��J���D�oؗ^u��Pݤ��
=�����;�v���e�����F(�\�HH�rT��������������.8�}��K�Np�q	��cM��y.��g�\�ſ�����T���ʑ�Yz5�;�}Ӄ�֥Z�O���Qܼ+��K��;E��Z~^R.�Ǧ�k�G��*u���7� �E�H�������R��͌��	�GH����G9������b�	~꧁�����@"81ϑ��Li/Ͼ�ޅ?9`�"�f�uơ�{�[Hj�m����+�	+]%�Y[)چo�Q�0�]�9�G�	���Q��z4:.���Cj�}`	���A4�m��Y'����h.]���/��tN�Ҿ�i,Pg�IW%C_�E%�>9�Ҝg�:4��;�ZBxCؓ�2�{�;�����E�K�k�tVl�U���m]�i�5���s�?�p�����p�R��p=��I8/%NK��H|�	��lWa/��W����`��~±:�T{�7�+�������3��G=��W�Ў&L������G����{�fQ��QmV��T��j�S��mZb���!�R>[�.A���B|�����:�Q����ٞ�ݙ���4(������ۑ�M���uQ!��u���{�\nH��pTr��L��SNW;�dI���G#6�lo]�8��u0��[�����h�Y�=���G\�^̮�o����d�1�����wi�k��O\&��#���@ .��B-�y�%���	_��qi�����V�9Dĳ�j9Bb1@7��sE�u9�n;�1�,\eTT������;���Cr�n��n���f�A�a��A�K��;���uֺw�s��O��gg]ĺ��o����P.��v93�V�">��4�-��YO��yNσ}NWd��n$r0M�c��O0&䨫'z�>'�J�:��X�N-��������qf=���
�8kK�;��+�X����e/\���?�)P=cwg6�⇲q�_Zr�'���C�ں������z�a������]#�8�&�4��#�&��0@���'��t���b!N��j�e�ŹUj2^��|�����aџ7�]7��E���!����Z�9$$Vz��y�Ĺ�Eш������Jt��T�_.����5�g�Ϟ�z���>(��{?�Q��@� f�)k͒$-,=�E�w3��PFH�L�����}���&|p���g��2og��`f�,�u��j�:K�L�SR,ۘ~��u7�2���+풘J<r���R�O=.�s�*��io�cL�z�L6���9������^�0�;x�n�g�V�4�~�mO��|A�t�W����<�ʎ���)Wmv�����(M�����D�IS\���kH>��%�d�zud�o�"���N���f���s(���y�k�V���Ɓ]��ڿ'5�A�}P�Ukp8��3����7�2�l2b������e��>��o-�e��%}�8���	DHQ�H���P��m�����������������w���6��������ӝ&-�^������i���w#��|���b���ێh�Bʡ~��fK��<��z��'c��!U;��� �� 8-)ė�������'������F�u�f�+�*ύ�t�^�Ҡ�.��������8<�m���ώ2w��K��7NRW�z�����!��劇���$e���jC�jì���0��g��H��3H'�l��x�廽�cDe��B-j�����H�w�S�Wc���I	I� ���!�w�#����[�
=�Os9�<?����#]�G�O���7EA_v�2��)h�it�sџ��s�Q���<۴(//?k�kᅇ?�����	;�w�9�9�-�F�Tf(�����7�7���IVt���98<�^O�*��/�u=8Wt= �����\���-�o�;tW��\׮��Y;r*:e��i�p�|��L�h�A�ߨq�	bH
�� Xo��l�]2�Ii�y��k��C"?���5�K����r��^C��I1�O�����Z3�s'&��6���R&�\�����6D��eխD�y|&�aݩ��T9�$z?�k(�3�Q�����g�D�p�P9&rXm���<���$�p��A`=d3a���\��MnO��z�i���2�?�ŃO�
�=�����2�l~��,uYQ=�
�����\pԟKAW�-[��QQNH}���^y>{�
��'���#|$�����'�5��f������:�o��.a�?��}ΐ;jĶ'^��w>��uk��9�<������5�g	}�9v�p�!�w~lW��Ra�xo�ac⾛��_~�U�ed�.��2$�(����� x/Q�g�hׅ�o�#|X@zW��j[�]HDEAp
<�?�t�3��B�뿉��'�����J�~e��x�A�g���v*Μ��Pv����Ț�)7j���i?\�W�Đ��k�G�79Ŀp�B�ˎ��Y�ҹ�N5հ6�t��ʍ]u+E���h��.j�轰j�pX4Œ�0���ޑ���Uח#@I@��D`mV^3:8�M�q���g/��ƟVD���������"��uS�y�u�f	xd<b�����fw�\QW��vokOchL�"-UEs��Y�Ё>0�"gZNj�
���L����6K/�7]�CU{��u��m�.'�O�	~�Ѩ1�|���R0�hlN��u�ou�ģ��
�2�������r|%.s�2I �|��X�6!���^���]��c:�vjS�xP�E��c"~<�\�H$�# �4�.�4E�m�1��I}�=#Enu.e�H�����ZMwNLK��(�����' j:�B�@�ggI,1 q��P�km�����#DC��{1L�����
5�x�9������W��B�8��㓓|��jM���T
1�$�E#6�ė�3��qBY9{ױDԒ�i���:������:.NL$�	�_���_�)�ᓄ����WM�
:*�&I��0J��w� ��k/�i�����s�'d&����w3��N�\�fX�l�z�"gİe�թ7���$���Ҕ&��1��l�Y�}o��͂��2y��?�s����%:$n��ҐZg����Q�ӕ:�bm����<���s�Mo��R�x���!Mo�+_vv;��̗I��tЯ6���f�$�n�V �sz�ҾV<�ü��uH�k��H�)��h���j����b[:Q#{�L��/s�]n��<[�Yv�*��ʓr������^t����,?~šZhr=3k&d�&���/�K4I��TA�u���N�����ڮ�T\]l�Ѥ�r�;�I����	IW����x�K���~X��4�+Z5������9	��6_uߵqTg�9�3}9X6��)G��r���C�z��v���j��i�KqS5��b������[�q�����u��ğ���UR��8����T��='1�4>���.qpp �h�>�s�9 6�H��m�n��H���n�ph<<��~�)���S76�_�Q�P��d9�K���{���4�Nf$�}ceR��eɝH�p��@Y'sO~���o-AE�ϜH㞴�@��d�BF>)�<s��m�z��(�F���j9 ��j7��I��/��8���^�����D��5-����qX)��N��w���i�7�����u*�tmz�,qv<�1�Pܩ=vgX^
����n<YVA���*�����Å<�&�ƒ���Ho��]�ׅ��d��9/�����zVp�	�.U��vُ�cޥ�i�׿�/QYy�n�Y��5�g���$��Cj&�>�O��ͣEr�������������2=�K������Tj�K��O�]9�ce	N�Ջ n<�y�"��%��Ϡ,�
M|�d#Y�2��~9Egp��E݇��]52

Z[˔��:��їͫ�Ň���1�}��#�7G�p�Yb�E�]��\}����tTV������J44��V?���}���{�Y��w!Ede����v8���/1r��m�`������NM��L�`ec#�����N;8P�̗��s=��罸{��4�4>1�/(=rS�(p��t+g��R��W�[R��Q<рG}M23-K�k̋�{
uI��N8��%ku��]�(�Ξȫ��ӫu'Nו�!���'&<fX&�d�� �f-1���݇7�����
�����=�C���VV�sG�)��"���#���SJmF%?뿬u�x��0� ��K��qi�Fӫ����>�]jpg�4�)q���x�}��q^SCBevqQ˵>-���7ulGU�6s�ց�بř�n�):�v���iEi�^�!���v�)��B�X,����q���4�\��	5'�V���qM�rN�z~�r���XX���hD_�;���5*�H�8���Fෙ5	L	N�S�E�_/��"����G��WۅW�#Т�lojJ)"��U�Z�5J�;S�d�E�.�����h>�i��D�Klf�����%�+�A��$:Ъf硣��OϥIr=6]�ĄC��Sa��چ&����>���<�!u:#9ĿV�9�u ��@�ȴ3�hC?�����8�Q�iR��S�W��S&,w��1M���G��3�r�����5$pZ��<����/a�ř��h4�EȬ��!�IG���+�Y��!���4z����>���?y͂��gukz�ߥ�r<�)�����޻Yu����
�<�7���L���cC�<�t+ÝE�I'�ǉ=�)Y#~��l���ʚ�ȑα�M�ՙ�[,e/��@L�fn�a�����L$�5u�+�ƞ��>Z�T+<hB�դ"�������4�U-e�<8�I)�m,�q����� �eY�}Ŏ��B0�@v���o�I"��� ar�q;�R���F?�mN�N��$@bj��&T�w]��q�cV6+�2�g���9��''���	R�3;Xe#y<`?��^n��3��$+���m��sm�K?�H>�>{�j�L,��zW��&ڭ^3c����b�Ҙ_'����b�e��$Q� �K��I��oK]�J]O�����g��w֟rC��p�X$
!^s��;��8��u��������2E�h�C�F��y��<�5e.b��C�c���ύl?ݘ�~���~w'LE\��ǻ��t��]��������]gzΜ�7� E��G������Ⱥ��T��6�M[]vg�S¿P[��#<E޿s��^��'�����*Z��.������|u�wD�'+'�a���S
e��k��ͭ�m�MY��ڥ����7��_�{���B�wP��l��zs�����0���ն��Ŏ`�V�A��%��kU� h����G�É��e&�)#@ݝ�P��%F���6��������{V��a&RfLhAV\�ov�9`z�c��%�����2ʑ�bj8=f����y�#u�,kP�j��ᚂ��]�$�6��	�Z� � i7"P��W��u��Dk
��i.	�؝Z�� ���Kp��?N6cl�V����4 �ʯ��?랁��֪�X|P�F��)��v +bvl��^ˁ�<ӫ��R0BRSS�~
M�����c�cY����2�(�r{�O{���s���Xa���R8��,��D�N�C�ȧ���T�	��መW���0W��
g��w�A�A�zok������2]�J�A%Ƽ�凞�E���(��)n�3��"�q��/}U/�?
u���#$���es��0[�T����%�-�L�z��;�����c��{����<���LS2:�z���"Ge�╼�(�Rw�O��)�k>��}�;Ī��ѩ��IPT�K��vm�F��&?�7nCMT쓏N�~�z`j�af�l�V���{�t�K�.Y�4�./������$���C������?d��l6q���z���E��#��d�v����U�9�G����=�m���G]+L6Y�_����� �݋�i�n����8Z��ܢ�~��8�p�$U�@|iD�R[X��df7�j(i�^@�Vcܔ��n��s 5��xv��r�ӗ��G��R"��,���!n�']��w�Vwҁ��s�R�6�]���${���}v%\<��lAy�|~���y�/�i>�>AK�$����M�'�tK���]��>�?	�Z�2��_Ү|�7��CCm���a��VY{8̘�LE�6��Ɓ�|.J/1��Sv��r���-NE�D(��]�0�4m?��K�F��i���kt�x>��O9=���i{���9��8��VRgvMz♂�I͸�������;��'�&z�ݿ������a�,F���Hn����4���3��V��$�h(7�@w��DE��wE7M�:��C��ު���{� �.���r����Ȩ�䘷e6*[y��]7-�d�>����)y�۝���J��~�|��$�:���um�*pfE��4S�q鿻��yͶ�*�;�h�_Կ�BR�+4���YM$w���!# �E#�g�o7[\�7�u�wCR�[]M>@m�Iɋ㡮���c�)�������ʘ������J&|�ӑ�����-���g���<���+��tAטs����#�6�j���w�\�Z���2p_{
�U�)o�>�猠S���A��݈�7���P�#R�����sy��Q/}�)��qr-�+㧁>M�c4�pu��;f��$����4?'o�*uN~�Goz�4^!s��|K���g��WdYY9`,[e/�&�WD`��ҰNX� ! 9����mtD�#��i��@���+��H ���Ջu���n�����(hiK%��L�<h�Wn����25k�+��KL�^qM#m�vb׀���;��[�E�뗫[�y��?�[��?�Wؽ�D�'�H�:PO���R�ū�K{���$�8�u���/|�����s�ΖD��Q�tfRU6a�@y o͗r��RU���8{%8p�W}dh�f�\�d�DK!d鴩uOD�a!-ŦlX���4����kڈ;��$�3�6�j��b���GO<�-�:��޿��L��ŉ�q��x�9�1�rԝM��.=e��2Ji�4zb�(2i�5�d�o���(��	�T��6޳���3ks��+���P@�4�<b����ifP�T�<Y��ХhfK$!�����{�uKQ88�N
*�D�x��X���Pr
�g�R#|m�Ƌ�\� l���[ͣ��6nӚ�H���z��u����(���u"甁_]G��~��)�ʪnD�/��M��o,�?�M�k23���Y#�k������1�{%�,kG�|�c���,�_	�)3�Ku��ٿ�<4l[י�k�"7u�����[���6P��),��E,{�k����&�������t��p٧�i�p�Ա����#[�g�% ?h��FG�e�zHB�O��F���fQ��ԏ�ruȩ� Ā#�%Z��2��������8����V�V�-�Âڒ�o����sܠ��{A!!�||�tN���e�n6-��hm��S����mҜ������g�~�+�Bnoo�C���''��z�����FO�|�����ǅ��JA��
��3�ȑ�1P^�a��0��Y�^K�Wl�T���g��[uI�Wǩ�����������s�{F�'N/��Ŕp��DQ�8:?�I������wT�#D�����"f䱎U�5ǫ˵ �Sr,����T��t~C�sᣣ�e�����W̆��~RF#%�G֔�B����P�Ӈ��V�q�&l�W���R��'�D�N��az	)
n>>>�~�R�mlOJ]��j�w)vH�TD���Z����csss)���t�d)�+BEL�H͌	L���������s=v7�Z4]���Q��PAƵ�rL�18��ʗ�J`P����~Ȳ��I�%�Gh6i@t�0�r���\l6���",��[�T��S�%JPkV�K5�c	��.��$E�3��=�"k��9\�m)t(�cZ�Uq�y��O��`2�Z��;_� �����u��&��u�٨�)!��2��4�p���e�$��҂�K�Ҩ�%֊�u)��~[�񔳄�����`����� ��;��L�]DEY��ڔ�p�	��̣���3��)�n툫�'˱�������|*`
ނD0�:�X��'J���'�L�<߳�k.�hUh��ϛ�BbR��D��~i�du�O�����R�X3�ɚv1��q��R�_��$�œه�R(�qծ4��j�� �p�`�6�)�1g�y�S��JX'�TjMҝe9�>;���
�85(�[y�t*ߓSPX�8B.iC�������4���C�Qحf�Y�L�ez0����?hP빊��h�z�^� rY�����p�fGh�v>pW�H��
�;PD��T^�7q�
�[�'Tb�!�|#��d��3��XT��)��]�*�XG{;_���l�izS�6y��r�xI��Ť1ĩ�x=���g�bU����`�� d[m@�͍�:����,Ai�"�p!=b���6.�L�\!2]=N%pB�d�4?��ɴ��*�|GWx܃������R�~���^!e�����Cg��"J��W�mc��(���`�Տ?�]7;����F?w�?�I��}�Ok����?�
M'�o
���Tď<�k~,��\/�� ���f��	J�@�J��Wpv�e\�#ˈ��5��;E.x���<I�],�H���2�ɄM��>��W�:�����f�1�r�{��V���$��{�Y�6l�J�={���'ax�/�+}3>�'e�)��Q����4�;�`pӮ�]ΌTL]\���a�w���A_tK6��b�Q��0ҨBM��l� ���^5��RTvAA�Am;i����H�����)�+�ß��I nh�%Z�,M�7И�>p�H7��M�bas�
��]��(�T���Iuu<q�.�s���)UPP�f<9�S=��*y��ا��ȡ2�,�R'�&�-?��V�C�f{{��ܼ�X��}%�ګ��V?��Y�:0ΞH	��¤R���zP�j�`��lc¼V¼�Ͻ%�����9#K!�1o��"�-����}p��>!��r1^��܇(?���e����I�܊h�qc�"�U�S�+C�g�s����}q�')�������qf��@���]�(�_�]$�g����Q�8�|��sdO��O�O�v�ա'▔��z��� �'��FC�� ��(OPP�QVt��By����{:���j����f,sv���̺�Dj/�9�<y f��~�����Tړ�i�� P�U8H~��Z#�_����wfyY�d;_��_H�{Q2��f����d1�X$)6�)��	&�������<���p�����K�k�>lYq�g�֒�,O�~iRr�e��ժ� �Ȃ�f��Et'x\�>�����c��F&�)�fe ��}�_���F����i����o�j���ǒSco�ڳ���ĦJ�֬����G,�C@�7r(��9"ZH}��Q�$ �O3u$��"{c���,h}H����N�0S3��{��eJ���{A�H:|)�~�3����<�(�Ӡ�>wb�֝X��;.R��Z��ߏ�i�Sk��K��D������K��Lx,˕��u�r��#������^^S�k�B�"l��D�{��I���M�M��H�P���E"ì��Fb��߭�f��Xz8�-S඲����-���3�Zkǩ�����k@kH����pc�В^����}���n� d*e���T��χLۇ�G���D���
��w���R���} �nk��z6R����fV��T��P��nb�-��6���V=����im4A�2��V�l���a)9HAX[�p<��D�#�#��p'B.���QE�F��L�@�4�KS���13�إ 1[��"e�2���HK"AAɱ�k��aK��P��}�*��J(?�U;��8���YV� 2�{���a3�ww/(jM�[���k����55_-Q���^>3��cE�(\-�û�u'��Kƒ��6]r�AR��c�T�TH}k4�^�#�~�9�6���i���vXX-�n\��Y`�F�ѝ;򶵵��%��3����ÊDw�� ���D�~���/8�Y_��g&�G�|L\J*ǝ�$��|�iYT��<a����H{uu����/-���]iP-D�C`	\=\��缸v�xؿM�c�ל���#3�S��I__�����������°�����60���Ay}��V�A�3�y-an�c�\�����H�=�����OH)*�V>Z�%r
fo*Sr,gŇ�:p%�2�֤Ԩ0	�agt�1����;�/�f��&3�0(0l$�9sA���RgS�5&�*Ebr� �%i�KYb-��8Ui�����ivK�,#X�؏x���W*v3�x�P����/��Nd�6g�}��^�}X�;���A �F�?$��)��u��`�D"�'ܽ 4�D1>:��tS#j����|����.`�1�7؜pJ
�j3�C9x5�Co�9��m@ԁx%C�c+��4��5�����%��U��p��h�wG�?�-��gzU񛪹re�]���1�1ѱ��U��K�8uc܎�]��/�V`N�-����^�>���vm���5w��+��c��^p��0��6��h,pV7Tm��C������2�T�k�MKXLJ�J��[_'$���zO�O�I��n�џ׮t�LemA��$Rz]
���$� Lن��9TTt��X���0�KlU2����v��&�v��Ơ����*`܆|T�ε�����E5e_�]�X0�C���Is����j[i�e�z��dw7�������Jbu��Z8�f�[���
9Aܲs�G�:k��G~�X�L�G�Pu�6u����]�t�p��ꓓ�2���'v�U5�nskk���Q�q�z��Ic
�lz�|�1�/�W�׹X�>s� UVM��.p�8�45'R��mn����+o~~~3�/T�o�����������wa--��46�46��PK� � �_�z�a�<���n�������e_s��T����I�U(l�p���ڼ>����HM�{�o?��K�YtV�z�4P��ӊ�J�~k^>`��up��-���:}�ܺ7� I@!�Ճzɨp�F�dA�_�y~Y�x�H9�b����S���&u�⛌%`t~@iT��@6��-��ZgY��>{�|r�f��I�O��f �;��z��e��VXui|�b;��	i�J�Fo�S7'<�!���K�q���_V�����.�yi/�s�@����Ҟϲ�F/!F$qsk氵 ���f ����	j]��宸6ٚ��3�0g:���w��/5��5�	;��C��ӯ,�����E�x�V���,��=���y��o� �mT��G�qM#T��W�Q|
���@/�;�f�*����y�uٺ�������/֏��#ji��M�xI9c�h2�.��?��75:��m�����@6�V j�r��$�O%�uM���p���.en�e�DөV"PDb�Td�����&1z}w=�{^6�-�^:wd�Ѳ@F6n-P6K1�R��'q��qME�S�t�c�K��jU�U+k3��)@�'���++��?�̱4�e`qm(�I���*WSӕ��en�h�X,oF �Мc�4���	��H���Ŀ�������.�Ȕ��2ĤЯ�X��$���W�=��΅����,�ױ��]��OӘg�,%M�I��l�PV!��JH3G��Zm=��ɲ���?�����Q�%_y^v^�9><�*���XO[�����6u�>�rR�v�����D&�z��|���\����v�Z��1�ģp|*:*��r"�+��s���G\�p�����D�P�'��l\~�+�녒�S��5�^�2��.�J>dqy�`T���jU��B���sM���L�(u���Q<����US�V�N��40��Tbĕ�X��Nǌl�:+ӧ��������"�qmm�u:�`&��v���5B">		 � �F(�E0w"e�c���,,��� gF)�se_])R���W��m͑��فv�^�2;6��� �*�ی�2��'n7?�.�g����)��<�������Ϗs����{��Y� ��t$qK��>��֒12b�����/�����	��ͺ�RWh�^�V����d�~��IA'g�Z��j�D��4���/�4���x6��n������s��N웡�#W.�|J����D|�JT�O5���{�CG�#�e�� �ĺ�������ej���j+��Dpg�9i�.��͘��G��{�Lv�Zn�:k�Qj����;�|�݀���s�����aS��yjt��i�������l]�q��cZnr�e��~����-;g�#��5�{���!q��{n���te�Q�y9U�W��'g��e���=��II�cM����F̹#al���JB4����)��D9����n��LqE[���"D�0W�4���/e(Ưe@��������w��6/��&)�܆xi ����	��ǍŖ��c�c�qWw�r���r.�����ؔ���S�8���Z"p`Ie�ӆ��v�ݦ�~?�Q�@�2٦ؠZ@R���XJ�+FcP���Z�V}EC�]�t�:�1����'�.�N�]��J((��@㸾�[�4��0G����=j"+"��oi�t��П�/7ى
��l\�P��Q���b�S�b�� ���w�@��dW�Uܲ�Eq�YնF��#:<���/(8�3�L\�b/����- ��@ÙrU�yw�I1�g)� Yyy���a������8���[ ;5OC�M�eN��WgǛ��U�"�.^Tg�L�tV)�A�÷�ί��k.d�;�f���A�-�WS"� j5���"KK6�EL�W�����=�"��\<A)�R��C4}9���<G~�b�7����xP8}s��j�z�͢��,��KI�W��!��ӳ)���a�t� ���1��DP�^��J�U�P��`�|o�.�Cղ����`$�XОP��E�F��3$tf��+)d����i V����/�h1�a���	m���_)�a�Q
�D���Ka��x2^aYA�G�"2����k��t��Ӵ$Rm����2y=w����
sM��]<\U��<c3�ceHg#y��U��J�?nQ&�y�1%[�������m��ӯ#OIk�P�L	cd���W
 }�̥4dT:��]�H�̻�5���P�?���"�1$^o�x��#+�@j?m-6m�6��o���ʓ�O#�ի7�f�)��i� \��uI-�뾜OJF�\���� ZiBX�3\�L�7�� �ؒ���:��QH|fV~.K\/ו�[�t��P[�P|j5$����yEne����[-B�R�9&�!ΊǼc2����	Ǆ��WՎr4K:��Ð��ɔ��?6���6� 2xH+o�o:���x)��i֟���cl	~����l��Q_����z@��b����g�q��H�_����{�����B�3/�1jސ�|�B]��&�x���T��=�FN1Rs�N8 aa���Od��|rEX���Aest=#�t��k|qc�D�m`��N�%�%gZ�۩�\�
6b'�&��1�GMSc����Ni8se�,�L�
:� ���"%&T;y��̃�<^�/��#�#�79�yeC.�1�)�iF�]l�.#Q���u��]�DRmlm�^�αOH��ډ{�q���v��/W����S|��B8ɲ��ݬ '�~�?�;j}J�`���+�$/��q6g����/����}���'�/fL6v0[!�}Hl7Y��K���V$�[0R�`k����As�&`X��~
�
�G�a�IL)?A HF��� �&aFr�: �N.�\5�m�i�	��5U�㓗�Z!�ɥC�]��&�$a���Q�*7�H���oу~p6+�]����&��s��A�?���X�;���ʧ8/�61���[nv2���*���������(�x��=&h����1�3+����E�*୓�L~oCX��<���3���jǚ�sGl!8�B�~wpz\dē���e�h�-5fr���(D�A�;�2Y >�K��N���BV	(A��ڂ�n���8��,�^��b�Iu2;7w�w ��j(�s��=�����M�z��b;O�;�ڰ�OPPm5aZ6T�߂<v�I$9�y��U,�-�(�h�6P�T�S�� b܄xW���5����?ӥԒ	Dl�n���/1LH��[�Р�ʁ�^��IR��\�F�3��D�lT㥕�����X��U�XY\�����O�!)��I�m�R�f�AO?��Iz d�ʵ�g�j���f��h-NI~�#��	��մ���:���=aϳ��WE�@%���;Ԝb\��m2�2�.9�7j��ܲ��27ౣ���eR.�X��΄q	��֛�J��̧qQ9���M��{~�$s����^��h���Q37*�vZ��m�e,Ζ[|��c����O,��7�$�'֋uV��X��<d�M�:[q|����0��=���7;���.�-��=Ч�⾺��z㜧�"[������ۜ:F�n��;#�1�:���e�<�G'cr��O.\%���T
zI��l����,68c�U�]fy�l�v��7��9^�Jo�X���LAN+TzO�ah(����{�l�&99�G�%�{<�`���5�B*�{��rppZ���˽��ڠކ�vX�RC0��jg�G,�U��0�B9�Q�8�ү������i��U�1S2ˤu�3.�����e.(�����C�96\�E*Ե
�Qh������ ������_��[��A�Hw�!dG��ip���i-�ӣڮ���O�J�C�N$`��=��p~��OWU�`�]UTF�XL�1�ߪT��4	�H0@��F�ʤ����3�
�6���J�����-�xl���u%�~B�^9�"��Ҳ���m�(��M��}c)��CI?y-"T�J�Q��� -�3�ԴG�� 2w���������B��d`��^S٬=�
�� E����	���0UdK�\bu�J�;����5]`����ˋ<�?���ZjV���h����8��xt�v8�&͉��0����W��#��L��w,=m
j�
tLˑA�j�R�٘�i�O5f��\�F�!֖O��i|k��Vv���G��e4�,���@ݗ۠��������[,���72,}�L��N�#Z-5��䜩��ѝ�ͨ��;O��PX���������[��B��'��^�I���B�j13��?.�:93�_�G���Wg��T�9?�V�<:��ڍJ?fS3 ���=Rx�a��׮ё����K� `zh>�<P��_Z����
�d%�O�]��|�[�M�2F�� �6W�����{����D�:k�2%�r�j9|������Ұ��+INyh�{���Q������}U�{��O[�����C�${��Ę�Jc%��윜t��4&S��ϔؘ�ˤ�j[H�$#(��ʰ�?ZIQ;�����t��8-�4�-���T0���J�)����D ��j<�K��OPV&�|a����0����.�1�7R�$JY3��(l���1�b�L�=��BŹQ�Y�6$��m:��ܥJ6�m4�]��*�bpOg��:ut�NL�Ձ��M�gϻ ���t�@]�kKj`q�v��w4�J��	�᩿lb�. ��#g����8��>Rt�%�.�x��[,���A#�ε����f�H ��RQ�g+���>@8sSF�фN�&�H��[��Яh��x@2])�M����wb���B�*9M����d�*�^iP��!!��VU���LwO�e�G"<�')N�H��_1640�
�{�U�[4�=gW�v5�i��)JIe|p�M��"��I����*�VW����1�?�t���O=��J*r�)G����o��=�]MZ�QM��'�3�H����G��UHB`���o޸ڨ_C_�5�:��c�%��uRc�4m����o�ȗ�a����(`�Oi`��qR���r�ܲ
eC��6J�{����צ1�e�Qo���Oo2�Ν�L�9�6l~9[�ͧ�K��dp��+E�cAE�F�NJ�
�3O��z�B���D�p�ٿ�L��,�쟯.MH�ҭ��s��"�0K��Z ��D[]�84�1�Ȍ[v댲�6�o[�~�䉿�h�\���\��x&���ߠV����%E	�,ƿ<֚�Z�? ּ��&��������h��)�֡tr'��9�F(Gs/�����:��JJ�{�E��<��V��_H{��5���')�L4�G���#���9K����I��p���Z[d��6���B|CA�ݚE:ֽя;�^ Yȗsm���QĞ!`���i_�wE~x�'���#���'�����ߙ���&Ȝ;A�3\8c8b�HB�N��?r��ro�Ы̉�зU��T�-�#��YAUN�ߜI'��+֍\R1�����;襖�px��:>MN�tx�A����`���z��gF?�O�BS[96�X��:C<Kƕ+L���(-�88YT�����9�C�!dp�Se�}�R�����3i�������P���ꧣ�D�a��u�?"\^�u���	���I��Q��D�t����,��?��>����^�gs��:����D��[��,d�Z:[��
��9%�S��?^�Y �$^H�C1P�.g=���6a�ȳku��ca!��7e����F.�N뺞ݭ�Ą|ߤ�_1�j�ޘ�[2%�5����9"�r^bGxL�C���J�����?(�g����t�ѨzbjI�Ah��ƿ`L��O���ĔĔS\L ¯�|2��=�*�{�,����W���'�}k���;;�PUZs���~U��	�s�#���Q0�`C"���L50�h�Ӕ�n�>t�Mz�JZ��LJ���a����qj�� �U�0[֎Ј��s.�S�b���dZ��;����v���X���D���C�;���X��7��Fo	��s�)�qt�c��!h�K�Qbq�_K��*E�ԭ�k!�agG�0���2������T|�D��Y�����p��HV��V[�ꂘ�hpm(�ŋED]����8߶9`��w��`���!9P���qt�K����%Og@���/�;0�-��a�	;�	M8�"�γ��C���($M�d���� �@F�do���2���>�p��g���;��Ő%&�RYPY���Ʀo֦	�T�0:Ed�F����!"^���C�Y�
���(�y|��,���yy|?��Y�������̍C�QA
��(���F*C�2h�ź��b������x9�x:�	
h���X��{�Wa�b�np��o�s���9���g��R��V�Y�@����$ o��yo~�d�����v�7JK'�`��aT��zD�Yy��*��=tlmnJ-�*�����*��ւ�:���E6��ػ1F~wD�Hܪ�z(%J�G�d�1x�'ІqL��7,�(�����8K�6���t���]y+�%�d��A�X�'Y�� nZ��~��,6o�7��$0Ÿ,'�KiN��p�]v�-��$��E�i@�֢�4�U��"I�F������Hz� ĭa-���G!ō'�Y�+v��.p�c���Q��<�l�l6��@�壐�E`I���q�����O/����h�3X���4F�QA�4�O���͑|6~�1����#�8�:�X�R��� �����l�$��;��f�*tFDFjU�%���@C4@�3�y�����0�QV>�]>�	L�`w� آZWw��ʪT�#\����\����,�� �a�|nz������{�>�#�Em1�E�L&C��3���:Ó��dD�2-�)�c�&��mm�dE�V��͗)�]��%�%��2y�G�X �-�����G��e]t�&7m����Z'�ե��6E��y�Ga{�Z=�4�)�1o�0Yk
�)���2��G���u�t8�Oy�s���{��w���������7o� �R���9�O>ju'<�C�p�Fh�O�p�� "5��Z�1�q�Gi����E��� I G`�\pԓ� �é�~:�Qk��ɳ\�}��;�$��H�	b�8�~�|v�����ZK�=�b�e�p�# 
�њ:����X}Ⱦ�ғ5�4W�ώHr�i�����Cb�h�:�G��Zm��0yN�[���e-�f�Tc���Y�y��O�#�$b�3�f߫@�;{!���N�"}�)����ծfks���u��7�󜺪8::���{QUy����e�=+A�Y4/pe�eCDe��tc&:�r\O�A���/.�mY���xbp���� ��`<�* ���<�xWr4�`h�Ԑ�9�ѧ��O����>�ѿ2)������������ ��C���4��Q�@v��K4���|����Κ��4�d�~��h�sB�ߏC �5@r� ��j*���y��I����:M�z��gy.�@P�>�,ȵ� ��c����>��]>����m���	��X!�h��(���o"=k�OTl�����d�p��i��|�K���tJn,g7���o}�W^~�˗.�g=Q!�^�-��o��|��?���o��9���V��Bd4���6����	Ya�!D�"gyi���z�E��BL�S&�1U]K�I��ސ�$�H�(C^ B+����+�N�qx���A1
a��csc����^�t\R;��A��R�N�E��"�lf(�������e[��d<����q���,	1b����U�ך��uVV�YZX@��3O���>�����?�:�ӭ}9sQFF����������~�����%B��ӊ��C��}�Q��<�!\]s�ƍO&8E�������x��x���y�&�N��d������w���۷��ߓF��U�����+N�M�B�k]��v��������9<3�(-3@L񓱓�Ov��E�#R>�'��Z��h�����.��ug��=�
�O��O�]��/�,��>���:�}%wX��E��i~�JO��\�	���ONr=r��ߧ^k�oIe1F&�1���`�����}ƣ)��ʂ��_'�O`Tr��t���{�/��H�{�����	�ޥK,--Rd-&�)�Vι�[������
�/] �,��XRF@4dy�/�~��}�u����=�Ʉ�U����Mسg�(Z,//������ӪB�H���HƊ��ܿ�&��(1H��|�9� ��*Yh��t���>����Xp.,,������
�Z���Pʰ�����
�N���d
41�h#����F��ј�tL��!��h4��sy���i/�4�{��y��}�s��������sKUV�ߡPh�q���<��������<z���݁QqxxHp�����/8�`�auu�+�/�����o�_��i��GC��}�Ϳ�7|�{���?�9�ѐ��QV��Ђ�ײ���D dD�d�EOP�^����>w���O��?�o�1���Ed�B�{lK�������t��{�(ѫ���d=��h�^2��/"�O�_�b<�i�=;�{L/���:E�f�6$,�����s7w�ӎ������\~���3�N	8�3�&	m'�|J�̽�4�)��N�˗.���H�*����^�KW���������x��	�^�Z�FyQJ���o��������98:d8�n��Q�G�H�U������*���~��g6���}�.���M�P�$E�aN0�y��7yp��{;�}��.����}�?Vp�)�����77X\X��JBX\Y��s��u�&�Ν���J�/�#x��4��jˠ���w���۷����>��Ro	�e�����2�^�j2�h���x�[����ɟ�	��,��Oz�fY�R��t�p8���/�?��w�3w?�GU��P�k�8�q||����Q��y�iz���91�O['J&���q㹛��?�#����/<���YKp�WVX]Y��{2��TU)��9=��P��O>-�'�G���l��(�j>A#����
b41�D0@V�C��y����2���!��� ڔ�g��p�?�xJ(n6N�����1��񧇝�#$D��E"+m��@�P�%f��5:�(F�ՐG���^>=�,I�t~,���Dk�V�M�-1ˈƤ�>� �kQ�BzM���,d'�&��̢s�	G�QF�FK�w���QI��lJ�?��&	��(��p�;J�f��<'��,˸x�7n���_d}}�N�'�@�����
�NK*'By�@+M�'�H]�G҂���+�h�ZK�ӡ�s���t�*/��<_��Wy�嗹q��g��p�<�/������p�s�8w�<.�gc}���b41����V�Մ�Dڛŏ�b46��Z-�E�g�?�7n��+���/|�[7oq��E6678�y�s�q��E�_<���g�βvf���*�ˊ�d�����{�x4�,�Ԅ��h#���I�ۥӑN(F[��������sϱ�y��ݖxfS#�:�p�!2�LM&hki�:2�UYS�S�	�ZxrOb�.���bz�����N�]�������+��������ĭ[�qf}k�)���V+ǘ��ḋ��p���p(����ǒH)V���ON�>/8��ZRT�������C����!o��Sv��y�{��MD^ǦV$c��F���C2�����xr��1��(U��U�5$>:fR�D��Y�/5�T|o�A���|�3,AɎ� 1#6%���FJdK�+6��.�����X>͈�g�����5�t'AKٌU��(eD[UH�N]��`�F�fE����gT���,�XZ^��r�v�3kk\�z�kׯ�y�,���Z-�\b����(p�1�L��2]��y���1�{ʪd4Q�>x�<�z2׭���]��KKl�=��W�u��o\g}]\��v�N�G�ӥ����uYX���I7�̠�'c&�	��b��+�J�'���<����[`qq��W�r��n\�ƥK����`aa�VѢ�i��]����iwh�[tڝ�^V����kF�	!zꪢ�<�(+8[:�6h���
7�����k�=�E�ף�[�L2�Q��d�Y�L���� j�v��wJUVTuE9�2�?Rpj��<��5C����K/����
�������m�[���s��e�ݎ\�0b��|�)~�Ƒ�$	H�ߴ	�\r�i�Q
�e�����kP�h��T왋$@�JD:�t��
��?b�Ѫ�V���g�è.*��X���ê.Ju0���blb[�Pt�:��ū�z
�j�"�6Ju	�*'�1v�+��z>)Aj�ĭc�����AFHYÐ���e�d�V�Q�r���c�(2�n�ULFp
E�1:�=��!p��ۄK|R�?5��J* �Nb�����._��+��4��J�d�HkM�0�q�#/2�769�[���:�ђ_�|��sb\!UJ�����,���=w��_z��/ܤ�[D) JI��K�y�6+Y�r���%�^��͛7�|�
�,�)��B���`cs�˗/s��u�66R|S�ؽ��R��'����\�p�7np��E��M�:R�Ϻ>ETP;O�e,-�p��X�y�ʹ,)�*�����l�R�$u�^��-��u��7n�����Ғ�����P�ǽ?#�"D��S��E�l��I�h��j���~�,��>�""�d�>y#�\
 �YtI�%�1�-��xѴ�|�(�O�S�p�-8��gD
-4.12T:db}>s�����G��q�8���>N�˳��V��	��ܓ1X�̷*٣V\��Ry�
b�
�SqP�(�.f����?��y��Z����#�/]D��1u�a��6�C���V>�D�Ѵ�#��#��$��z~�h(̍�\��1Y�����iw(��x���1���&)��g2�0�9�3���v;��i�[豴��,Մ���ʌ���$+��n������&y�SM+�����tBUW���#n_�s�iT}�?�U�8�<׮]aumu���i(�H�第����ϳ��E�բ*K����＠�(��"F����O&x"��]���a���K�Z�����!0�L�v���,K�Wk\嘌'L�S��1ӲJ��O9::����x@]y�1t�V�WXZZT��{�S��<}"���b:�rp���o�M���h��{;;l��PN��R�*{�|"z�ǞbMʳf;Ĺt��y�v�%H������|^�;�&�^��"��Ȕ�#h�J#蚠#Q�xpZ���0	}fg��!��'��1��%�p�>��� �W��� :R�g����i���Dj�������kklK4N��QZ���(�ȸ�6���`��է�'E[� �4
�C�r�@�j0�=Ay.����Nwi�_��t����?��O#�4y�����GC��;�������#���pp��pBY9��0V�Z��b͹D�z\0���b�t:VWW��ؤ�n�g<�0���c&�)�tJY��'SF������`0`<��2���Y�X��$I��RD�k�=Ν;���"�ʲ�,	5�ѐr\R���=�����L+���\�hL��,�YZY��nau�B�O�#�*<M	��v�\��hT���d���?<��p���=��9>:��p���}��#��!�O�D2e��i�	7M�Ȟ%vzڕ�"�y6�������-���g4�]���x4���G�y�}ܿ�p<��=�9�5d&O7�7DT��{�*�A����<�(B�#g��A$����D E��8-n��Q��o�����]�=^{��� �Iڽnc#�?f�x�Q��N`�蘲}��( ����y��k��=�Fd��#B0:�����'���`RffR���Ӭ:�|�����53��̷H ih���dh�_���s0A���b�"jR��ĂN���GTmA���>�LTkQ��Iu�3�/p%�L�4��Ȋ��jTRW��#�\4ܠ]O���w�M�e<���������fww���=z�Σ�CVe95�����K��*-��e-�T7��(:�+˫l�o��L	4����>����h��ߟ	��#9>�K�Z����E�7李#��e�muX__�St�]�x0������=93MFL&��1�~����w���LJ����6���fV���Ӏ�ӳ���W���V�9�fZN88<`wo�G��y��!;ۏ���a���}�GG��s��ݔ��k��X�MO�O^�F3��������o��}�{��曼��;���;���;����?��yp���D6��|����i�i,�+R����s���ދ)����aC��)I���5_�Ոl���M AX�*	�H��h<!z��tDi�
���쒽(C'��lI��3�)p��4N�C��pޝ0���x�<�{�I�_�8�;�3��N��I�����B��L�f8FQ�B2���t�ň�Q7s����	���@AJ�ފ�B��Roȹ!bY�9FQ"�����~S#2�Q?m��ʔC��tz��C�E$@�x��qT��W3*)��>h<J������s2�}�St0��*��[d:�0��G��Je���$O����`�t2��^~gTx%nG�\�|IH]W8�R�aI��uB��JFSq�s�w���>��p|t���UU���'��(�QbA�,ߔx����I�2�"�+���8W�e9��rSP�%�<��Ç<z����v�w���cgw���O�j��*2�VN�N:�X37u�6%U����&��jZ2��q���r��d!{�Nƌ}��	e9%V5��6�Va)Z�"C�G�FC��HO�߇yz�5�;yI)����~�]���o�g�������|�/�����?�_��ͷ��-~��F}*/��	��x�d�}<=y�"*@7���3�uBS�-�KlP\S*Hۡ�d�Ր��8ǔ�Bt!%�M�ۓ�AIV�hȒ��(�>�Xʔ˴G2�7�O�@H�C0��$Y5�ZT�}5�t��]�ҧ�-C��b��d��i��<��M�܈���F�:�*]�)A�Xd*��bz-��� {� ���g��Z�*���3A�}J�c�_;J�|@����v%��R�|$��Fܡ�C�F��A��}Q�1����3�J#8PN�u�=����/����A��>5*#z��h�:J(I9NI��O6�?t�+:�2���P������������t�'�{\RN���I���pxp�p0�rr�(���LK3�i��NK���A��OQ�~�SU%��Ѥ�`4d40���zZ#�(���K��cA�1ɳ0��8��Y��r^NK��)��QϊJ���d41��9>�31���ג�� ֞��P�F�&U;@� CߓkP*b���t����������'�
H���@p�u��	��E�j��M�37�j����T�YI2�T[�wL���8�8::��>������>���/��O~����}~��<���Dk��iZ�f	���P%��'b\��'���<Z���2�ϭ�uv���k����a*j��ĨQơ0��p����c�Ƽ��}���L�5�d�:Xh�/��/.Sq��f;�D�&ĈK��"���3�:HȐ�$6���7��zr*5���������HCi�ZJZ���ojH'�'_�U�~��dq����5��uD#kE='PS=�'��{�qC��3�|�iC�29��<���e�i���N	 �W�/��qNTc�w���|g���GD�����U�����B�ݍ���6�u���cdJ�0�
I������j+%V�w��)G��1L���J;���"h���H�Rc3b��(�A��p��]>��<zDL�0��W��xĴ�3�#Xkh�Z,.,��vYY[�(Zd�E[C�5U�(]%�$�x�CI��vx��t:]���w��e{{�~�d2b<S�� �$�� 4�:�Yz�+K+l�;O��!�3b���`�x8|�p��U%u2�b���ڠFcvw���>�'�Y9JL��&�;}V�)�7e9%��6�i���-�y��2��4P�����]P�p���������8�ߧ*K�ՄjZ2�L�O�V�(3M9���<����$�a�n�"-N����h2�Q�[ x/PU�x_˂7�$ ^�m��	�g�hp��4�T"��X�R��(Z9׮^�k_}�/~���/�kg_��&� ,55by�^����jM�����o��ÿ���ͷ�9<�l�3�:` ���>1raI�Gt���N�f��1�O�$�����2�B�!5��?Y���$5�J�|���5z��_�'�澜�N����w�c���Ok��3�Sa��xj~��5g==�
i����5�#t{}�,s�,kK�O܆'H�+�i�����nE�2�~����u�4�0���Y�O~�YԬ�����2!y�hu�\�|���"y;Ǖ��s[lnlpfc��<Ih*�P��UňsJBp��v�%��h���Q��!g:���Cj��V���U666�p�</��2ׯ_�����)(֓:i��|�y��j�Zs��=�~p�_��l��������%�m�>��c�Xk�t:l�;���v��n��ҥK�z����,����EA�Xk�:P�, 8:8��������>���G�vvw8�quM���k��}�!���q���ј�����ι�XYYN�A��?U�GR#��̂�ܿw�����(���c���R�9�� �>���Zcb��Edb%5J�V �����<�Nѧ�m��)��A6��֛c�A\�Ef�z�
_���|��\��D'�h_bU��:m�H4�IP1L��&�����Yegw���yĿ���wqt<Ae-B̨�C[a��(y��R����8$&E��I�~:Sk�����_�R���i������԰��\A���0������U�������^O�) )'W���v���OBɤ�JPxҩ�3��(����ro�e�lS��G��`�����t��T�O��>z�4��Y����t�?��mV��3����\X$+Z�G}����t�tZ�qT��Sg�.#FQ ����ǌ�Sƃ>y��++�w�9:>�FA��J��ޙ3gX\\�̙5._�ĥK���ڤ�롐x�~�>o)6k,�@]�loo���޹��ɔ�h���{{{�#�_M��֨�f]�bª�v�lllp��VWW�z����(
l��{�O��Q��k����w8<8���3O���e0P���d�g5@�O	ΕUVVW�L�("yQ���L�ݑxi���(ިfŋ�$�K RO+���LG�s(c�������ÃC̯+8�u�#F'`$A5�����>����>j��uJP�Xp�h+ҷ�9^%�"�S�H�i�\����_�ʋ\��B'7(�1�D���`R\��sL 3��:���]e��o����������mst<F�|ȩ]Z�x�\a�Z��$ �,�գ1� �I�bMⳓ�����-��"Uj؋���J[t+�~��)V����ѿ
�7<�!��԰�O!85%��x��eW#�����T�4ǥ�K��ѧTd�j�ۥ��/��,Wŧ��n=s	�I>������$>�r��&%������ӂ3|�hu��D^X��}�>�Nz`־&��L��5ڍ҆P;��t:m2�crMUyZ���d�����F	rOBG�
�@�h���L�ץ�]`ee���3,-���� (��Os�����3�NEH�ﳳ��5�W��y��5�$��F�,�YX豺����"y���,�����EA�e�ؕ�O!�R�Rͪ\���x�`��#u婪);;���M����\YYaaq�PUT���1��s��@	�'N�5U��h#��t�"Ҟ��fwo��>G����)��Y�
tLZRL��%P�OUʜUi��yҠ�XH�h�+�
���Ċ��E%9#Fυ[|����׿­���2
��]J� ��J8_(Q&�M�s��"����}�[�����*!�u�[Y�Q'�s��N*��H	�jX��N�� }�B�����5�+��j�I�W������,�ٰ+R��ӎ�����ף��}����ŗnz�"Ǟ��4�8w�i�͝脒;\�p'��̟���UR��Qs�b��5��OJ�œ�f���79���S?�1�G��S.��%q+�H�&�|����I��OZ��B�B$h�6�����i��4fn�Z3���iC��^����X�p�3w
�uӵ%J�L5!D����^ӒG�����N��������Ǣ(XY]cmy��b���2i&�ИJ2�6��2�r_C��U%�'ڭ6�q��h�p8����p�XL��Nk-�n���uV�VЙ&����V�aM��Ҭ:F�#��4�{�<Zk�L&S�����]��NR����HՄ��T�]@��}���.*H�ʺ*��J��4��#*8�n���6��ˊ���Ψ�Hp5��d<�������MNRir�`0�L|����Ҧ�);;�@����J.�q�>�~���J�>��B�y�V��֖�ta����>��x�����C���g�,����9>p��.���O���3)=���E�������1�Z�o�ʰ:�jG��������2�"�d#)IqV*e��ьu4��jس��ȴ��'�2�L�Ꚉ��@�F�c��YΫ�]��<��_���}jX��g�FI}G�Ғae�O>!b�Dp6�H����h�$��x��Jh-Z�����s.]�/xN��gQD�0�I.?!�^��!��)W" kM1s���ߓ�,�"-��? ��j.�C��
��N�r��S���w�L�n�����Q���r���h��\�r���"���Xy����M4D#^��{�I��#�����+B�p�S��V��d�Ç�L�)JYH�!�v���gVWYX�#Tu	t&��B����`G#�O�'C-Ir��'�F#����1��x*!���V��ٳgYZ^�h��N�����IfZ����ئҚ<����P�j��J�K[v��u�5��KUI�ư��g����!�4�*�Ҩ*AX��򈂨�&���U�R��(p���}���o"��ds��K��E�Y�p����)�)̲E��ASP��!D)�x��ԧ�eE�� iF
����+�<����u,�������_��7���;T�\U��<Je��L�F��"�2PM���ӊ�`r&㒝�>���������	A�ʱ*⫒��5n^��o�56W����6���o��Y�{%�Ԣ�������6?���y���p2m�C����S+�'��	5��	NE�F,K�y����h�h'�^����s7S�d�K\]b�>|p��|�I�~JfxHʏ����Z�'����ǐ����
Tb��kP��c���75})��՝�tClT�IA�(�Rk�(���s���q!e��'��N�GX�3��Up
0@����ի��m��)�le��Q�M��%�CG2���	�SU��UU��s&�)���g0�3��X��|�T�E�`em���U�1�%x'ªN�'A�x��M�t�zTZJ	���:��5�є���zN�S9�-3���iu�8����*&7dZ�U�s����8�N��ʉ5ƈ���T��ֆv�M]��Ӛ�x�����jZ	��2m(+G���������� �+��G�)�D$��*�m��	���*B�XJ�<���?8����ѯ�)�d~I?�Ȅ���#D�,&P��E�N��@wS:7�1<�Ĵ�AΫ��hI�v.�}���) Y&fq�k~�w~�/|�e���)�G��O9�*D�E1(���J+���O*�7[\ET5(��-��|po��{����p���>Q[�α
|U������.�G_���m0ȌAk���m*SjX�,Wa:��$7�:�wx��������8�FpI�wh+]1����P�]�=
N��w:���M��*Vw�Q�ףX��v��3�ll�K�|I�J�|L^k�5��L%�=��b<���O�/�0I08ͤ�g�L6W-������Y�e�|���>�f�={���-z=HL!$�C�dw�X))p&��,g��}�	I����>�;���=��fq��J|r��;4�*���o����%��
�n�,�R>�FG����Bɪn�Ri�e8��h��p�t<�%������jϬ����D�����c#:h�J�I�DS}�zSKF�!����H b�+���c��������"
E�g�d-���c�~:��Rj��*���L+���GL�	1J���@#��l�����ʙ3뒤���R�%���BQ!�p�Ai��cf]a@��"jW������{����'pR��&K[M�笮�r��ά���6�$�(MP�I��R�Jw�Q�jW3�L�|x�����#������<��5^}�E֗:��c2��2��d�Tj��AAf�uNYU��d|MP%ʴ�&g��;�w����{>���1�f��P�N�X_�����|�[��2��0
�
3�0̣dȟ
��E4J@�s˴��c���?�����ѭ��b7x�)�l�ʎ�v�ߓ�T�<��x��ѳ��<5���z��cd�r��ynݼ��/<���\�'��sv�O��yzʝ:���;�g?�޻���U�,;�%�B/
n{$�\�=*͍���gP��?���|�i+5"ٹ����n�˫���k_|����3����W�ل(h"g3!*�5��ɭ���}�~��7x���8����OhV⓫0>U�=
�C����$B�Ź��i��h� ��Y��X�OR��@�K7	%�I�~<���ˠ?��J���Hł]��,�,K���ԓ�OJ>%���5(�����p�p8x���(1"$��q�ٔ�,//KV�R�a�I�g��,
A�TJJ�ٻ>xƃ1��cFC��TQ���A��c���������ڪ`�F�V���)�D�ߠ5�C��2jq7ֱR
kII��������@���l�{�u{���r��.]�ąiw���-LV�}Mp�ډ��"��;��ie�rCn�S	j��Ǽ���}�=<��tZ���3��b��6y��r�:gW�	ՄV+�ʤ�_�)�P#���#��ǔ	*�(�aU���#޻�����y��6���Qy��9::b]���������?�]���)��G��C�j�I�h�✹|��XK4�:(�������׹}��c�nLADQU�0)��Iv$�|#8E_{ֻ���ylbA�Գ�?�L͚���Vwz���!x��6_�������]����s����x7�'L�oH<(�p�)yaV,�j'��8>>�Ν����g��'?���w�h��R3&�X��旄�$K<�ϪF�|����0��qRF��X3Jk����?����ܺu���C4Rԟj�T��l�*�^�_P�է��y��Ϸ��-�����}���&#��g��J|�*|�+�ũ)9Hb�O�O@��[�4k��O�P���A$ ��A�Ϣ"��=n>'>.E�e�(�%����F#��$ˋ�=��#�H#�N�M��3x�yoՌ��a���!��>x��8�8:<b� ���L��X���CQ��v��ܗFᘧ��g.`��ٜE�RB�֒I����LJ�j�t:�V`JjdQb�����t��:,-��� 0��`�
���EHe�2�_��� t�+����D�Ч���)'3�oĊ�1!�ϴ���;7=�˚b�E����ŋ/����._����2AV`J-�����'�V'�9=�s��(����x�����y��!ñXw�	�,.rik����x��yz���Kr�qHiG�r�)����cDa�T}:-�R%�3�x����G�������c���Q�"Tή�p��y������K��T2�"(�A	XwS��N��.�UD�1�S0���w��7��!w�?d0�d-����,���gs�{*�X�ABN��t<"�f1�h�ɱ
N����yO�=o�5�H�re'淚5[[>��ӌR^���x��W���~�o��78sfm�N�3�:uZ�*���(	21��dH����x��������7~Ƀ��Ρ�᜘��<ƴN�&�-Ty��\=N�g}ڹ`���<B(M�N�������3nܸA�U=�Ut	*�0$�FgR���ͩ�t[��ZY�p<�����W�w��}&�qJj�.�9dOۗO��>Dx�D��,�v~�?�R�Ƞg��^)��Lֺ�3���h����<��5G5U�q��D �1FjW3�Lpu��3%�D9Kp�,�j�<O}.֞���P��No�ذЄf�>��u%ͤ��Ę��N���:���V�zM�Zm�O%���������:�?&��u��މp�ˌ2��d���jZ���fd��O"�Ep�(�ɔ���x�P�G�Vq�Ǩ0i��g�����$�h潑>%8��~��d:�3*���=&3F��f�bK�Q6D�t�܏TS����͛7��W��K/����[d��t�C�A:ٛ(�C ���!}��$�yі����ux��w�śo������'l�<��K�]�ά�G_�/\���b?��c�,N�pg%&u@��5��q9���P��~�����=���?���><ƶ:x[�ܔ�sn}��\����׸u~7�p�"S)ӧ��,�*�1
\��)�%ڂ�;��}�����Gܾ����eJ�M�����OL�q�(Q+�V�Ԝ)�\�PYR^NV��>6���OuQM���)�Rtr#s�J��lZTQb�i�d:��'M>F��5>FQ�L�^���%o��c�"LEpvx������?��o���*���ȔP!
�]T�੪���(��IU�\�W��d���~�U������c>| �f�C�ж'HU�M��GX�3�9�g�':�����f���^s�b
�Dx�y��gu}M�]F'��!��{On3L�Sd�e��Ab�	Q�#�����w��7������2�N%�<s��S��yz���YwͱP_�_�jj�@2'����=Ǯ|cL��J��:
���԰�jf���;���e�!DlܳH\.A��d���#Ƈ0_)c���P<���$�)A_SJ,2c$aM>uJp>���74���4�4h��	X�d���F�L���̾W~�|���>8���8S��^o�K��I���6H�Y��5��1ڀ�#Z��_�ފ�#J��q�u��R
B*gL����d"^�L'��Yl���J�SR���c�r2Q�2��蜴k~|BpE�
�W��2_|�5�����ٍ-:�UU��b��rr�ct�zN3�Z�����*MVdX����~������;��B�B��֙e���Ë7�rfa��tDk������"���.(&��n�6!-�G�G�}�����y��6����V�`r�%�M�:��W/��_���oP�	T�=AiL(ͯ��S	�C���`�"ڜ�k���h�����ܹ��A����N��+|E(z/Q�\���Yl�?W9Ɠ�,ކ� ��J��X�A.2�̈́!i�(�i�F�	>���5�wL x��Q�&M�4��d2��O 3��h�A���9����V��_{����|���eqk�H�M�X�U>rxx��q8�3.K|�X^^@ac�����G���˩��t�@��uj$<Ϩf���&-��8)m�1q�9R�j��j�&͡V�*����0ư��H�ۡ��dy�J�+��aq�#/r��.�K���zt[�Y6qc���9�`0��o}�o~�/��w��dZ��e��v��q��l��S�'	φ;S�3T-ʖn.�)Y6��Ts9gN�#D��.��R��L�X����P�-h��"JTS4)�����*�(��0k�%�w��!F=y��.��%�,z��d�~�x��ٟ��9�Ǟ~]�TƔ�3/EB�BS�%��e������O�*<J2�g��ɻ�5R�Q�6�l�R�\c�9�G�Y�-�/eY�\��0�'�bD$u�E���kkkt�]|b�>Dlfx�ŗy镗��˟�#V�B�p�%P��~w��j'�EG�R�Z:����եo�1��NJF�1�>���p@9�B
8�Z-�_����2&����D%��
ҙDE�-Q�5-r��
k��xo X��)��C>|��^�p:!*���A�u[�YY�����YZD�H��X#Q:[H�M,Dq�7n�T�*
�%ǃ!���?d2�Q�S�9�2�ܴh�J��|}��/_����͛\�~�+�/s��yΜYca��R�=Ӳ�.4L_��b�X"1��B��l�瓻6J�Q�������k�R,,�������k�x���x�7�s��5.]����
�^��&� %"��0ta8�����un��W.s��ڭ6�J��5)�$�d2��������po��h�d<�Yn�)�#�҆I)M��h��vA+�)�m�"����n��v;��]:���v�v�C�#��jQt:�:m�EA�ݡ�n�n�g;-���n�*Z����S��E�#G����m�"��j��4�-r�<'�
�VF��!�,��3���0�F.�𕧬�Tu�d8a<��1Z"H�k��d����}��o�����ŭS�[S3f$�6�Q�N��!Ǫ]uT_-����Cpi�+��A�Kqw����.��`E�kq+ZR�[)�~��#y�$���ٙ7�ξ��r�����Z��	b8�����2ױK�J����y�1�Jl�п�� ;k����_R�<���H��O�����hH�"�r�X=`��$0�N"V{�UpAX�V��#����l��s��9	\��S�M!{���RnDF �tPD�d��3��\���9��At�y���BZ�$78}�2�{��;CqF��"�=����S��7D�(!;��[�7���Aav,"H-
{�"x�O\�J�5�o�XS(�0�Ff0�e�����ֶ������`k+�d�?�Ɖ��:ӎ�߫ص�2*$2��vy���z�d���Yr!�(��X桏O����x#��
&�[�^u;L��{ĴD�W:x�9}����Bdyq-�
[͢W�P�Q��oaN5��i��R_���{	7E�uv;^��:��>�3��#o��f��ɩ��M9�d8��^W�|_�(�4G7S��\d��E�ˊ�p}`3�8�j�����f3 Q��/��isou���G�9��v?��L�o���1�^�ԢzWm�-uw:���_�|�G�ceL�yƘׂ�����Zҷ�� v׾O�2���I2/H1gw�c;i̒�Q��2
2M��&�ڦ�e�03l�B�S�䍆�-_��C	��4B��C8=X�<VM]�r��m�7���. ��%JA-}+f�,�K.�'�
cCU*�	�5Aڈ�:Z���qlD��h8ԉ(l�s-�3��}z�yr�o�۔�f�<#o �#f��WW*�B�Dkі��P�6�X���CtK�yX7vM��{Q�eQ�w�LZ:��W�h1��GF�Q���M��Yn�ԩ��:��uSl�/��m�;Dm�д\ˏ�J��j]/@�9���c�ܞ9 wF3�g�s�gl�ѳ��� �z6����Z��Zӧq�_y��	��7�VL�~�~�7���� b<��W�.O��H���P)�dD�� �	b�ص��p�2�N���NH�Jv%�׈7���;��v]Ss���8�T����oe������k~ �K��������"ܝ�9��7#b�[.B���m�ыߎ�z��o&2� �ixpT� ���jd����2l�(
�8�ȍ��K.�Kn���"HX�bȄ5z!Vя�mڃEL�/��\|Z��{0���k�k�����n��P"�>����!@ݝ���b�g`��b'P�����Ϟ~l~��/u�Wճ�G~v٦~뼹��g�?az��:ӫ3�މxe�Q�W���>���NY�>��(�4���1��I�u��U���Z���D)��;�JDt���g���ķηBGH�O�H͋lY0gX��$�+[�V��bt�.��DH�~�!�wڍ�ˤi��aL�(���z�������b��V0��my��������(�¿�������i����蛲L[��$&}�G���F6�K��������s�T������'km�>Z�8�� r����nL?x}��f�����~ ,�E鑸\E7k����F����Bӈ��d�U��[D�&��������$���e��^��h������a���� �j�|v��WЊ{�*����
G'tP����m��� %U�����xs�5E��۹������ß���j�������k@��yL���8Id5c���yL>�v4��bl��qw=���#����M]_/�96L�Lʥ��֐3���W��&{{rn�0Z�o>m5ݿ���?OO�\��sї덬�#��7�^��΂���Q!,��95`l!�ŭ��_�(X޼[_9tyc.���G��]�(�gǥe�v?`����?k�0`M�\@�$"���ׁ�r����E㟾�j� ��FA�إ�^X7�����?���>G=�y�B;�m9j��AA�j�6K��jɀt%��z[? ��Ĺ�
����푩�46KUF~2�¢yx6S5����&�i�A���������R���F�f7_)㗔˴��o+�%��
�,e��YP�s�k�+F.߷h�΂F��QJf_�Q˦h!D�jQs�����a��"`4���UQ;]MG�+��2�c��j�q�����:ԁ)��p����-Y��[�l.�1�\ɐ'k�OV��[�Rw6F|F��s"1�����pg�QM�\����`�(���E�%�n�״�Я��dq
��s{��9]��ש��zC���\VʑMn*~U��T����8���+������}o��9^�����f��kMy��Bh�i):�+�k��`�C��.���X]&b�������,�L��)���I|���r���歠"�؊#�Y>�Φ�`#uU	#ݓ�����la{�ф��ؖ���u|+Ň&	ʞ �f��P�ڭ�3��n��i�p�`�_��#k�M���3�����;i1�?jBt��P�{�����������ڨ�+b���Y�����c��W�X���O�O�"��p�T�LlcU
vp�j���M��X�i讦֜���'����OHuN�8d���2w�VУ�A�l~�ZH�>�ՒO�C]�m�����k���>�
Cٽ`f�g�>�=Cz��?#��tr�-{u��;-��]N2c.{ާX!^`���f�]�nې�P�qf��6���8ދ�i�VK�3����9h�'Y������6g�C��dn���:5�M�sh��e�Z�Z|t��H�\JL���;:&�}��4}M���~&Pl�f�!�J�k��N��73`W���%Q��IÃ�P�8�2BxR��(To�	��'�p�����N<yyGIM�Nl`)喭N��1s&��Ʈ�]����'ZN�#��z�<A;nN��t,��й�=�.��F�F#����[tB�2������W������>�H^'E���zrآ�/T\��ń�=�I^0� d�S�t�^��䆓��R���[�h��\��G*��46!���J�b޻�|�klҰ��i��2X�^j��Mv"#C�Ũ\��cti}�"q���S6���T�iT��x��V���j�z������C���o۽���i8ĵ,�l�A��+�c�Ѯ_��
GW�\����j���/�ƍ8��l�~��gH�¸*˔e�0��_�/����Q�[>~���{�$�T��q�PR�)PӍ��Φ�}�C!��Ǿ� ��ҡ����#d?��Ó5)��P�7!��N9dT�b��#9���"�����4�Z,�<��6<�h��l��/b��qO��"�"D��ŸT�;��
��Zց�4+���s��}aߴ��Q�~���8h�'ߦem�7�����	�\,�w{f����Ы�j<9�	��!���9��^�qu�����-�ڻ� �\�%j ��9�����A�����`|�EF���Z]�6�1�硓;��D���A�L��g����s�D��e߽ 8�7�"���N3}΍��s]T���
w63����<��.���/��(�n�m����v�Ý/�yiV�n��}�����(&�wt�]��G,R1��"�ʧ���	%Iv�9�d�$���ri�|�����~WV
�Ev�"v��`h�`��%[�^4#�:��-奐%����/�f[Fx�drK|Fw�]D��A�p�g�O����|�l����#z7dH՗�3��ɔ5���y�+�6���T����U�tp�t�l^��bo�6���I&L�K6��Y�8Q�� ����2�Pb�f��6H��>��� ��ܩ�����+ޮ�CS��g
�u�u���1�J�:�r�?�Sy����b�c��/h�F��l��p��P���K����i#_��[����n��	1YL8��s9���SY�f�H��O����Y����Xn�|��Z��É�����W����2%�F�ˆ����s=r�i�h�:�����ƈo�뻧yw��	W�������nd"�Y[����Jݰ̦��P%1��[[�A��A�.3t�.6O!�p��8�ޠ�u��Q�ϧ4��X�ʻ��/�Q� )��
3(�|,��}�wgﶶ|���WJ����O�L�eyL����1�?ѿ�j1���ML�qq���l�9iDt���"��?쿿����p?��kBΛ�������d��5޻܏3r2���W���<#������+a��u�
7q�s�.'?t��3�s�}���a*���i1;����:�Zi6�ό���*���g�|�n����t�g
YY�0��&~��VF���Rn���.Ҍ�Ua�0=�(�������5��-���XS�k�v� �����_D��B����o ��ј�AE�B��W�%�b��f��KZrj��hOY���>��vu64v�8��}����Bߜh!��t8��݈@�lIɒf";,����(N���*4���oB����xk8�8`{Qﾶ>(M��g�P�w�4l,�MH�&ҫ��{5O0,��Ϭ�o��J�؞׿'q�.��g+H���$΁�!j����.6�p�|�C/8��$��3�)����>g7�r@�著hMm���*���
��at�g��)EHE�%����t3��haM1��2�0Q.��	�= �Ϋ1U�|�R��y/��MJ�3���d���w.B;a�t��â�G�}}B�W����	��ܑ8J�i:�ϊ��(�YS��38{������ܹ���{dv�aSǶ0��Z��ɨ�x$�N�%/�B��*آCH��4�r����5����K~��3�ÐfIu%ꭼ���E?�0�q�o���G�+)���wiՐ���A��rj��e�
�������a�/\B�S�h�C����(\�\������tVJGo��չM_�T�_�u��eZXYEx�d��

.���L,����
���[�İy�V��+�vw�ɩ��c�� #''��G'��q���B7	�8��$�:�mh��4)��%����E+-��է�SAi�ۚ��l� �{�s���yLL�ݛ�]>t4b�)t#7�w����
rO��e�9�Xо�`�^��}1 �z% /�Pv�����-`��*J}�J̘]ϊ��)����6�lS- �х4�$�)��T�3u5�qi&����9���X����I� N��Պ�'A��n �Ǝ��j�1�*8��O�^6�}��b��֤��&���1������U���W�����j=�G'�}&I|�I�lt,�<7����xS��8��rq�5�7����i�,���od����s���{u���s7'�DM����,��_��g��˵l��t
����n��ޢ��Q�`yۂ,��.,,#�q���#����	T�ç:�Ũ-�3Z���w�N�Ʋ�e6�_�X�֠װ�{���8��#�V�t�:\.P�^�! � -���mmmӆ�=cߟN���mtR��]L5"�?.AJJJ�ƫ�c��1op��gq}Y�zC߉d�R^?t=�vv]4\5<�NNN¹1E0b�ƪ��g���X\������K@~�HX/6�
�Aĉk��!P��c�L'� ��>US�"�-���zںVh;�����F��������eb_9���?�L�ϕS���*ǯr3L�R��y�N�W��Qu ��b�D����Fm�I�W�J�|ن]s{����M��k���:9�M&�
�]��:�-�s��ƹ���q�w���sx�Z>�88����/>Ӛ��C'���%2�8%��Ʊ{�yVJ�h�t�S�Ѭ�|r웝�9ޛA9ݏ�N: �b;�zF�|�\ǘ��L�hor!13P�*ݝͫ,�I����TFT t�K��H � 3�ک��ȅ{W�ǿ�`s�������s�|���`kr�5���+�(�Q)^�ʕ���ߗ�ɬ+����ɥR��5��d�d��Ň��k�93�)B3fS�p�����=8M!�����p���7��_;샍�(	� �|ڡ��߿m���f��d�[�+�:�0�!���������w�^����q�vL��r�N�s��XW���1/-�ji����g*��7��1m���u��y	�3����үT���6�-{��R$�x�rX_sC�So+�������'1I�-�o��l���q����`g��̦��+Lš��;�vS�����c�6��n_w.�z�Z���^�w��%v$�n|���ob��~C�2�T1����m�X��^�M:�o�#(��̱��q;�M�n��s(�{�嗰s�پ*GZ�zӌ���*i��Ҩ�+s��60�<ڔ�^�n~��e�-�Y��S'� �&.�F-A����8�N�����j�y�h�I%#`?ӂH���n���{Ҹ@,>N�i�z��<��QGo��(G|�������'���JBs��"R�f12��L��1(��5f迎��ϳ�ƶ6ia�ʀw��a�D��&܍��:a�����jE���MF6�ʒQܾ��D�l�����aO>�ƽE��z��lx�������z�PJ��~΃�Оש�T�t��ȅYD>2�΂;U�J��G�c����Ql��U���84����\V� ������<��]�1����Qe��p��v���h�8��X�ǜN�Sg7��P�ӑM�:��J�=�(�]Te��87+~�,v%n[M��,; ]EX�����Pa�0�@�JL���F��W��F(}��y|�&��:�j~��S^�4�vR�����jh�-�Y-u&��K�W�"y+��D_�.%?{�>������1|�8F�9�.��L��6Y����~�6�i�&����Rs7��,	O�Y���~.�u��NKL;?.9_���!w ��z�
�ՋR� ZB��j��e�=r����V�,ؙ.�W\�$��T�E\��ki�MJ���y7z5x䋝NW�X �k�L
�f깪u��;�:��|���'����?Ic�oL����ykߋ<�o+��_~�K��;��kD���;���,V��B�0W�b�|�슮���VK9�ï�ϟ��}<�`dH�z�s/�l��%c�m�n,X��_u�+ç(��%��1y�ay�1L �ɂ��=2ZSs @L���f]��aCR_X���y��Z�0�E�,�@)g#�Zb�Z���ͮ@��%(*0� 5��s�o��!�c�-F�'Pm2�y�<�_�/�C#g`����;Ğ�]XZ��i�'ɴ�+fU]O�A����`�`�j- 6�I�� �T��kb?�w��_b	�dE��ܠ#d�y&�U�"_�g�H�C�|��g�.2��{�O�M�{�2`}����J�::z'�.6��)]���2�r����4����ih��71�ɿwё��8��tz�c	�����zE�Ll�mb�
�ɚ�4�R����cIR�+�w5�+��aL+,�$R�Ҋ��H�T���CUjS[����ȹ�0�X����}��t��jM�{�15o�������v���&�EK�^{��3�7����i�%(�8��ewժθ���������F�i�;�[�s���{Z��C=;e:mYQ8\mό9*�[�-��؃��fz�� �[�_��ˋ�Z+�<#*˿fI�.3�D9�ߔ��=6������o��k������'@�}F��tЭ�p	P�5l'������3<��>�x!G�m3�PT5Gn�k��r�>Vݰ��	u�ׂ���25-����k?:O����T�R�ơ,���_\���������"�8l+U4��[��NK�ާ�pk"4�ߗX�̌3T!���uR�'��0�G���Rsq���V��|a����,��$<i���QR�r�]����
1�,��ݮ�o/UJtK���+���?\$���e:$|0W���cZ�ed�>��;�j��){�8��ZRX�c
,.|��O���(�F���O������*^smJf#�-�l3����O�2�Y!��Q��-��i�똇�5?�~U j�BsQ��k�M��
��)����ߠ�
������}��w���bEu��'47�:�8U�r�5�>��A���Ex�1���Z�b9��|Y������7�E����ȪOyJmz��5Y��09��ha���L_4�'Z���,�un� ��-���&L��ñ��l��1�?]ܹK�F�$VW�~��"0orR�ø9S�	�5���
N;�z��"�rsz䲙�u�r��ʱYY��M�s�P�g`�h�в���X9�=!�8�gS'��XSb=Ր
�j�Q1��;����J�����Jf�k����8�nO���������?�7��mo���<��=�"4(�*�v(�-0��,���{�k�ń���
����E`�>>���(��Q�44sb{�_�m�������_��X&s�qR�2�X@͎l;�\���ڇ;������Oѻ��O�����x�/�ҹ���}�ز��q�?��3��2X�ŞW�ƃ[!��<���9� �2��#-� �%��v�&�i��ȟ47+���.��
���n����Z����=�w>��q�ϛ���;����_�ǰj�ؿ/h(���2nPv$�o��$׋�{*�p����d���$�S��V��q�4�Fɖ�	��#��C�	5;0������>;W��۲x��pv��0%�1c���ّ�A}���3�e�&�6��w�k��?b(�1�A1�r�;m{-�Z��B��5T�ؘy{�6T�|��*ǆWΖ�%f�=։X��*	w� ���Pw4j_7���v�ꍲTr�8L�0[> &/(�:5�qx'_?�jt���`:���s7A�	z��VtЩ�iyi ?%ahH5��P\K"8�~Z<j�ط���B8�7�O�W�c�(λ�Z��RO(����q�/�R.�f�ϼ���!F(��ȶTڎ�H�r���:�H�.5�l_ �?�Uf�X�Mr�O~o�y[�D�+�&�Nz;�G���}m�o��z�ʝ���5�,e�_3LbU+�Y-�r��[�;_D���`�����^^�+++��69y�?OOGwo�::��lx<"�Lj3�%�"�T$�3l��z���~t�:8��ٝ�����	�}�s�*(��U�}�'�8����d�����/Q]���ǂ��x�W�nh�~/����8;o~{v>���"L��/f�GMU���9��m������wAOKy���6���/�����g��W��W�|O2�.��6wm�{&Ծ?�_����������.�;��(�*���v���lJ�܏r}�ioU��K]�z�WF����E�
��1���h�[�a�q7Kc�&}�m���W��;B�l7���6,��IM�p�7�s�y��׷���]{�j4^�=X�5& ���k�RC�_�	J<2�5#M`{�1�����c���汹bά�1/_nXn|ҡ��m��{}Ե7Li���i7% B��Ȓ^"���_XϾ�'����+n���t(+J�a��N)����|#���1���T���}[H+�*�gM���#Qk�����E�)+/��œ<F�Rk<J�ə����f��~��^;|��>Z.���Y|D�;H��IR�#�H$1�����Ђ�ˊ5)boc�����n��9�ӕ2xg�^���m��������.B��_/��ڧ]�,g�@Gt��6�$��[�e)���H��=Ck�)t���m��ƚ��s�I�;�ӟM�m�ay���<�8�J�n?���z�6tO�m�:�]��G�\�[���s<�|�H� �&Љ|���>�E~t����{��)/�	j�����ihf=�L9�o��>�yq>+x�l�=�7
߻��%��)d���r��/p����U7R8����-W�b;P٭׹Q�v�����J���Wtg�}���n�
��KR��(�^����r�j��YE�l�|I[;}�g��PT�3�6*,�,��݋L.>>k�U�Z�s�:7wv*�,~c�H�ٿ�+��}�HٔP��G3��( �\b%���E�{[��aU:��������8�b8BF�8םH+eќ��r�.����7g��Ǹ��SԦ~5�
�UԸ:Ԇ̐Ĳ�`Z�C5��<��W�s�N�^�������]��T�A���D7��;Ť��l��@�K���rӿ�c��������O�]��hٺ�[ԂE�^i���3'S�FD+���gg33M��f���:���D�ӻ��H�*��#j�O8	�L�)�،�Ǒ�<�_)�S�>���'̅�����b��~Ҍ-)a�zp�k���N񸸏O'�b�F��?v�Cͮ�0S�vm�b�%�:�+�F��!%���Qԅң�[�&�h�Ɉ���
�s���-�W�� ���(�F��,�PJ�Cf=���������7hi�(���{%�d%|0ˬ�["2UU�g�������y�]�xg��w�.�]�g(tN�W۷<t�.�hN���O�}y����#'|�����G$�e(ҩb$��gǢ�q���|�N�Q�}?��x���|�Bi���=��{�:����
����Z8?'L�;%.�iq'/��/ �B�{�����ѵ.����5b��`>b�e�;/1�u����oϰ��W.�y��Ј����v�����t1�UYm��h��Y~���	�R���w]V��:GeX�Ъ�#T���Hd^�-U��o�Wn���%�,�FQ"� �nW3��֔`�$���*ğ�{\k��Dk��J��K�]T)�~�;����D��(�W~Ջ�Q�5�[j�5ݽ(�W�j��ܭ�<z\ר�v��(~,%A�g~]JyM�x|����9l�@ SD�"�bK$èB�2���g	��t?� ��S�L��|Pv��[U���dp��-"�잻w��YV��f�`�v[%b�`V�E11�7P
1�+�H}��*q�`8�,xmp� �<�LE)xF�τb��p�G����FCD��~�B�8������Cf$J���xPs��e}LV��R�5�͗��S�+-��:R�L��������R�s&�c���N�A���(��4M+��e�|2�+����,�8(U��G,��̌Ƽ���W�"S��#�FK��X::i 7�Ɋ��m��l��Y~@�o�������>�	�Q��(�-9<��_�q5Ɠ+��
W��̱׮��d%	�Z�r.I|�م$q��t��}��{d�@�������ip��^e��2�ђ羁�b����ڋhg�R�0v`=� P[�&�N���^��ƁQ�G8j����9I-�k��M=(���r��
� �<f���aA�����/�+��Y�T�Q�j�e�+���Ȯ��H�����@���y{�[�����F�wit1��B�E�e���\q�� �����x�5��A0-=jUU,;�CClcf��l����#��ɯ�:����sF"2ۦmww����N�d~u�jX=���v&.��ao\JoD�X�U�n.5N�J��m%�J��*�%A �*����-W���%%����I�.V<�o4 ����`���1E�8AM^�n��>��5�*AK�e��A�AjIiu�J#\`��������B�7«{b��J�O'�gj���t,������y�$������O�ӤM���;��hX�U0���Nͬ�-Ş��L��x��H�P����݂+b
M���2��-^�A�1���Vk���<<[����o��,����=1C_���K���R3�}��C4>�����gy���%	��͸2�d/�\q�����^�@��e��(�~�\�z�����楷��O����偡K��K[#��X�9(O=���OYG*��Ĭ$�C�NE��p~*��vI��a-��j�Ӭ,/��s��\�G{�4�"d��6��z���$v}�Nm>��u��U1E:e��1��r�p$���q�%F}qade�b�Uim�0��Ks�I{��ܪ������^����.�_����d�`��7C>�2�"x�h�"�h��Ř�p�Sk6�:Sx���y��PѠq���c�F6VL� ë)��� ߼�l)�=�B㨐e�"I+J�TeY+��:ll���5���IK�;�L�i��\�_ϱ��KP�)�-G����aג� UT��Re<>̳�NJ$9�p� N���9P}��̊�`����J��bf�m��XY�.��V��V;��F�Ǳ!	���E"Ъ���ic!��@�Y0[B�GU6Z��x��\�������M���BM�VrS��Z��gdziTw�c�&ڗoG�ϔQ�^���SB�TM���.�\NI�.��:�߻�##�0"��T%Lñ�IP�21���Oi'�R��&B�l�Ш�P��t|���lA��)�/��ur�@Tͫ|Q,�H�E)�GĒ��+��T�b�5���E|giׁ��3�K�ms�K�h|�Rfv� U2�u���/�R0~-����a>� �X	�����C (��ω.a�a�mQ5v��BF�n�4�>8���ՙmF���"�&�o9#Į�*MWE��֧}��[�(���V�̢���c�Ɍ�*�^���䉇�s��q�$C��nת�(��ɼ�C���3ʫY�k���t���g���� ͢3)�U}s��%��w>���o�+�dsC�Mg��7B-�w�SO��T�5��򘄐I��!D� ���2�UM�d���1����Bh"�!*�i]L��黠��A4m�#V��b��	E�c�7�ÕI�}Bs��q�W�Ȫ�U�L'�������5��n��z�������fK�&�©�E��y���DW��;\��ף\vC�ُ��5��R�,	R1��<���Q�R�b����M�Xc%�0�ʊ{����u�/�}�ݮ
;��wE���ټ��_�\1�V��v�w�,��9�h��%�U��M��b
�O���^����c=-%�"�p��UN�_9���b(b���:����g�'�8�`���Vd�_=^H)iT]�Ѽ�b�ۧOX����Z��D �<��+���R�[[��"$�߂Y!7����T�v�sj�N�z�Q:k3ƶjk#y�B���`g�?/��l��b`�;pg�H޿P�C��ࢀ�yz�6��M��-ƅ�mM9�����٭�	R��o�5jʇ5?�k��!��B�B�9R�\�\���a������1|c���Ҵ�?�m�^�F_D���h�527G��8�`����p]g���@��x�b5�)�j)S�B���sH-}�:7����nw�i
j˶���;�E,%�G8���f���#�d��!Y��}W>� ݦ���i&Ջ%l�Iek��R��F�i��V�ʚ��su��v�\�~����g���OmF�§;v��T���	�~�����Z�C�d�<�I9�}���/���󖺗��w��j��l��D��e(5��S��[�+�@D1ن1c���0+a��2R�R���[Ŷ��$p�����>���J�y��$8K"���t���r��9��G�c7�?��^'[U�N�.����S�!��bƂ�P���W�"�\����f|X,�l��o�-c�رlm�u��A	1�9�p~��MTn9�s���8��(!e��W��V�>0�y������#��q��C(7��ʭ��٪ev���֍?THI#򮄴�h�̝&�H&�Д '�t�����jl��Z����#aH�q1kP>�6�B�G�)1*��Q��c�%�7Q��ZB<1	I�G�#����3�5��q�?TA����1$y�Q�D
���J����$|�b2��O"�L��$bEBt��%��a�yy{S��)�i=�@7���vI֦�z��J����|���A"%~�O�s�5�H�1.Z�ayjj��3:��JM��U�@K�*e����Z	#��,��x)�xA`ڹ�Cո���]���ӏRe.�q�O79׍(4Wd�a�����/	�{<M����BQ���Z�݂��i�X�m���2 *�z�iT�82࣓������E�ʰ?�r��Ii�hlvl��Ղ���%b�r��`��q��ZC��\������v���Xoa�J�8�z}����g�)U#�W�ҝf�����C���n1o��~�BD{�瓻�t����A�,U;�]����zO^<��U��0�C���s�g���J}�%H�פ��EUq�'�z,�u�y�R��0�۷�s@-蒸��/1>����z>2���-��Pd&LL~β�դ�wK(}*P��r�̲�T�/Ƣ��/�_ vl�X�ײ��qk�o�J�x�7u4I��=�LXm�3ݛ�q�b��?�w�[�jh�.l�"܄�?P��K��׭�\?}�5}p���%�ggr�)�)�u�m���V�i�pǊ����M���z��m�}۟Ql2D�7����RA�&�;�DqJ\����[��HQ[�AG�t�H�q{�ӷ�7Y��	�0�n��ӫI��;����T�?���V�~)�����FL?]y�� �y�ð>��n��\�qho���d���X"��3GH�j0b��)��-�"�h��w�t'��o�|û����:�L@e����}>�-���_>l��J���!)S�,��O�$Yl��	)�
@�~Ѓ��C4��ZveR�r0���bS�읜M�d34<{����8

��������a�xĪ�{.�u?a��%�t�Ϩ�%m����_������>��	Ͽ�$�v%������US{k��sN�<��uRz�j�'� �ݵ��齽�.�'���ԑ1Ov���
���b��Bޒ	57N��L[\�/q�$�1���9��>�{�#)���\�v�]����S:��;��W)�fs��a�����XitM�?��k�� 0ـwZN�d:�<v��du�g(�#���T�"��O���g���p��Ы��G��뜼������aN7@��n�eI	���K�{�=c�ӏW�O0��_�S�`�J��t,#	P�t|Wm����<ѷ�u�K��"}4���X��C5��j(ㇻ7in�2۩r�1W��L�=�![�mNM��Dy2ck���v�Z?s���"g�M��t�f]�>xKX~���\����B�H�^�p���v-�^�t��������-<KyXy�����B�5f{���oօ���Y�:0H�뚾�hD|P=�f=B:�/�Ts�]��qvr��:�6�^��Bt�32&$(�^`��J��^��1�����?�,�P�Oԗ'2�6:M��h�
�{�/9�����z��6���xz@������5<\�Nm�T��˙�a� J�q�Pb����y�JF�,Uֹ�R/[$B������T�i�V'Yf�m8i�� �{�p�]KF��,o)H�X_�*dJʠ�tDƧ]��h6Q��Qp�S"cKR���;f}yB� �H,X��5�%bXx�e���ᬹ��%pq�EN.|\�������ӿSy���h�w~�D��D1Z���b4d1���c��Ǵ�k��T�����k���R��B�AE��9V5\܍�m�$:���T�m��:�R84mt2�x6������c�2DA֛݅'ܭmL�m�#�V�z)w�PB_��E�VWU7Ɍ+�QBڻ���Y,K[Z������{�	����@��c��y�"�~��R������;a+��˃ʥb+�Y��w�V�	֩+�<&=���;DvHqS��)Ϯk_)_�r��?I�Vw��.K�����(���G�;Ŧ_<��}�9T�^�Qi!C_�����,@���*>}��$�A*�`F|��ϯ�/C�����L���0� ��HqZ�wⅹ��[4ɍ�����E��G��D�W�ܦ%��Q�=�������G=�|���"wD�[
�:��U�4*����D�su
\�G�+=���(5�JzpEW�C�y�W������������*��EtǟzEܾ��P,A�wd�c�����c\A�9aҒ Eҫ ���b�*?�|�>���a�/�=	���������!q��9���$�������x����Q��Ϛ_�L���ۃsX=Ow>�9�W�oM�n� ۋ���%�\I��N�??m�.M�������y�Rc����ل��N�Kl*;��GY��ur��Z�Z�[�)^�ٜ�>]A�)�T�o/J/ ?���߀po�V#��_|,��dA�`����D,�=�P)c�l���֟CI�59Ta>�`p�&�t?��9��	���l5��\��a*���]�_�񋅀;jt�N�Wo�|*��؛I�n���� ��2a����5P�\�%cd4_��R�I7fĀ�wT"
�XN�^I/���\5��,0�.��!`�EϮ��lT^z���#Q�={�g�pIo�߶������#�*��h�eBp����kp[��=8��$8$���.�!���]��_��_sΞ�=��5�O�LW��?w���2^�h��L0������t�J���?μM�3w��nW��m�R"�aL�PZ5��呬�_)	A//��/������8��0��l�)s��P�C�zmr x\���f?��j��������a�:�3�n`(2�R-��dx��Z+�m��)��������Z�i���J�
|�?T��F͢e��Ӥy���X8��;[��5q��|�B�ʀ?�����(C�����~#�HCvCȆ`ZE��W%�-�r���׏�0\2���Z@�{�x�*�ͧR�,{i֨(�RyҔsoC��ƭnڔ#�a\�|��a�]O�|���)� �x �Zs�=�܆�n2ڵ?���˿�X�w�A+in�}�GGǋ����������q�;j??�dʲ��	ݴ2�	��Є^]]Z�P�X^��=��A
[9�[yؕ�.O�h���'��;j���G��x�4;7{��`�NX��?����`V��w��[>2n�btDmk)z�p�c�B�h�r}*/�ݗxq��FT7�X�����EE�=}K��P�yTQ�`nn@�o�^�|�$Ľ��n����-yb�}��]�!�c�Փ >�Q۰��l��~H+���酯�A-J����8Á�>q�[����٤̿<������s�C�����!F\�ݦwh���y�����?��]���♕��yp�T���|�t��۰C6��;~��>�V����������]\��GofDEE�֚~6ݾ��ݝ%022ڸ%��󧾉���GH`��mR�@��=�Px���MjD��p�_��-��Mt%32�Q�<����H�a�,��:0�3˶e|6�_�q����M�+�o�L��g�^e��=�ŸeSk��?v������:�Ȝ�[����!��D�ک�����j�ЏLz�v�，��?K��&LI�k��N4��������pb �L�_o�|@�+�B��[\@P�}���T�%۵ob�7�;ȃ�-�i�L��I���@U/�;��ӵJR!k��r�?��n��pQ��V(i�儕C�g�!��(#fʴy�|�=�*d��^�Þ+ؽ����t�~�T?��c�]ܚz�
��c�!�V.�/7sk�*���nl�������U7]^M{��I������__�LA��ͰiF���� �4Yp��U�,=?5�9�t��/��������s�d��
GES`9�߱UJ�@�x-vM+ăI������&)Li�Z�����WҚ'�������1��j�2�}RV*a(-����X��#����Сn���A���{OB�lg�`>>���.!:��|�kp2΢Vɏ�o'��Q� ���������/~�	���Fn�P���^�����	Qs�B<�������1�C��N�˿�S���$^'+;��[�f����KFF�.Y��E��_�1o �`HR���=�g�!�-/�G�w3�Z�`>]�1�߆�v|�k��?�VD���!��f��l���v6�Q�w �MP^���t�Y�!{�q�� T˳Մ�D/I��F���i�(�GF����3!�>�E1#vl5O��v�s8�z^`�����u&�G�}�
���P��17.qp�bi�z�z����L�^J��)�)���y���w�82B�T�~�H���� ��G�;�R�5f��TȰ嘡^p�>P�����~,�hM�y��Dk|�/ۏ����'�3�6�W�o�����s(��\U@w�������URF:�NJ�:�"�|����rՔ7׶��	�,�^�F����3���K������i``�����?��"\=�:D�����2�Uf�I�<��h�	��~�D��;��'t�V��a�hF!�#fnȀD�nA�t����8a�%%��7��ɉ�ܨa�{�:�Z��w�m�21A�vTM�&'�T��Kj	v%�$�	�U��٤���3��#�j:���[���Q�ï�fW�4��&�SD�JMvm����,�,��0��5E����Z��w��>�i��948��şidYv˧R�H��T�գ���sMG�XʿŸ���̿k/���sK��d�� �3��x+�#�rA8�<�H�����@�B��K�?�����\��<xx�u���?t�����h�����C����*Uo{8�F�W*�Ԋ��'���a�2Շ�ƥ09j�頻�_b�E�������ͫr�=1	�y/g ���o0����G�X�s��8�&��)�zS
k�-�7P�f��+� 'e��AE�s�n;^?����nL�6��i��*I�5�l�y����`�Ɵ+��홃N%9����az���"��n����'S������ه���5�2�����,�������Q����J��r��o�*�3�??c{�:r?��c������-�`w���C�x�h���Kmmm�?����>eč���"V�y#�l��M�H�tR\��8�m�؅���<IT��>�;6)�x3��Vwe�[�_{K�5��1P�Q�� ��A髋|�Qq��Nk�B'�s#=��_�h�P��c
3(����TboҦ�ʺy���'r�[�T�iX�W2-
�+��:)�a6�ۅ�!O�{LXӹk�b���F�ȯ���_8W�muFq(w��vk�5G��)��2��*��xNՒ%��٬D��t�f-K$��nn^^��.�U�t{��ح��0�Q}~y�3�`��-�{��"��sG\P��ϋ/�F��YK�*����$z��,5W�c�6dNVۇ�?���^E��g�	x���r�����P�J����3��N�Vn
mLA�G8����!س:w��T��צ�L3�Nv�V<�:'�ͣv|?����C���H ��I��lh�96J:����0�#�U����*�T�O��<TJ�7B6�=�StY���Xe�;%�J{�&Ñ�_�����7�Jb�DRx�o8|ճ�y��ާ��B�"��K�g��72�ux,�����q�T����pi&�����;��Rk,����n>�B�H�p�gi���������R��Ue�5�W.�zA��V�1������m�~˲B�9�P)e1M.�C�=��R�_��#��X�z=���8�N�2���i���D�'a�K�9h����Es�!��o>9����d�D>���5�I�Cxn7aHIbj/+b3�dK�Y�H���V�mxGPȇ3�h�E�J�q��t��q�^_zV�,��4�q[�9��0��x�QK�@�N�!�~�oF��Ph�\��� �n�8T�h���$���v�y/ ��#~�cU�_ C^�N����0,e�hI̧n�	Ӡ�+!����v��G���?���H�I�Bmp�Q�8��Cǎ�*�dF�R�"��1W1��bu=��3�[J��ՕG1�'�3D%�L�Ƈ�!����)�q���˿���&eu��\�v�1U��wD�x��E�K@`��z�������K�ȓc�n�v/g�Gx��6�;t�J�WRڦP��ж��N�3*/�,+>q^:�*�(dĚ�d��VV�㔊�ÌocSyH�E�޳!���3=͙�Rɺ�]����(�Ӈ������M�ݥ�9W�Pp�.��Ñ��fa��棿g��!x�dY�!|�MGet�K9����`\��sn�/���U��"���y;�Z
�G����imy6����a�9C
}~�]X�R�C���R��۔d��1k�(,�%Sc��rɽD)���lcE7���l��8�J�6�������R�ՎjIhߘFy@e��,�q�!_Ӓ������=���S�P��h�y�j����ӫ�nd)?P�e���?��i�}~���H����9���M��i ��ge1!��ja�E��K�J��S3��$�xEK{Y0꡾�ڢ;Z,I^B�;�vK�k����!�f/�/�u�ߖo�(Vw_q� ��P(/8����!ܙ֙z��ޔ�"D����	1u	�₍E/���F�����N�������sy��F��r�Gx��|��s
E�>O*� ���sΧt��mA�?\M�(I��&�����rh�Pn	/����7bQ��Bͻ��E�
BN�,&��(�Zy�bp;	%	�4�7�_0!")=�8kX2�BF���b2���6<�;ʧw�Ŀj8e�&~
uLA&�>P�3�dk>S��B��B.�m?�Wg�rNa��9+��QP����%�G
Ċd������,�=��n�/:�	����$J�ڐ,C��i��訕qH�Gucl��،8�Iq���+��7*��UЬG}L�����Gm�7����$�x.:��
T�uI��ϗI;���H�F��A�;�qv�e�R�;R�Տ
��0K�k?t&���Ry����As�f<�!��Bpފx�s�qw@�ሹ9ӿzʕt�Ԕ:�{ZGh�\����Pz��ݩD
ew�.���&
A8�Ǌ)���&6{�Ɔ�� �`��q��n���΁�KB!���q����K�<����=�Ï�j9�������4���lÑ�B*��0���M2`&3.<���o�^%�Y�=$R%tR	�o�8�+�u\N] �1�{5���PR�l�oH�E�ϞJ���(��o��"��Ij� L"f���wpo�{�U�Qs��)�L2Q�QMe�^i�4�M�}�,�y�y�r�*f�G>�M_̫h��BKo�|ES���4��>�*}j�3�Z�Zˡ�yse��	�,���'�ҫ��W��w����D��pdeW�tߘ��dx�쾴z����p���7,v3�㪒��5y�GF9j�Z���brɋk0�0�w'��$��76��R�K���F��6m�k�Q��s@;�LZ.G�϶Ϛ<nP4r"ь�:����}7�7dN*J�6-����h?���u2	_=��ǂY�L@�����$��|ե+�b��:!nx�3�F���a�2� ��K��GŇ��1Q����E����L>�8"��A��oN9;ri!?Z *�γ��]ը�_�`X4(Wp�;�����b��-WH
�@���v��C�ON.������LM��b������:򇕓[PP�~�0�%|�`�	�&���@������n��ef��ѡ�: 1I�qb�~`�n/��}��m׌#�������Q�Z����4��L�a�C�����+Dw��q ,>+V`>_U!Kj���������>e��.�V����g�'>�+3K;|��R$	�3:�ЏIE@JlE�(��߿l�_#t!��i����V#:RI�X�}�"p܃b@}x>r�C���d:y
�8Jr.�����F�%e�f�6�s��2�aU��_��4asؐG'��N�t@AF~�r�Hb�Z��k�&��}��@�&d��d9{Pۿ�ZX\�pH-V\X5��"R�3S�+�;�b+C�����T)YV�����*�_I�LӸ���Qj�����XZ�0�E�2��������m�N�7�?�x����G�q�3}C0��ޑ|�e������r-'?C�����4�һSZ��<eeq9�A֡䭸�SZ�Ea����� 8�`i����#9�Oh���#Q[oDѼ��=���ȯ!�3�C{�A�/�@t��������f��g�gjL:g=��B�BC�*���E�w�����l�)�~�C@PZ���=٤����W��j� rMAzηD�&T��}Ӽ����l�(����D��S����!]���MBK[C�#^����HZ(�Jn^����-��Bn��1�i������A�~��_�j�����a�$q����nO��5z���6/��`Q����q��^[[@
^�թl���n�,#��Vi�����$ݚ$���9;W�Z����5Ϧ�9�vu������ٹ����R����T2Dm?1Ȇ��ǺYS�M<���uor����`o�;����PF���>@��9�J.l���h�<jr��o=LB��
�RV��4.,�P��͞O�~#�$�R䨾��*d!�M�#AH��n�&������"�T��XA� v�D�d�{� K{G�	p�����}Q6j��OLb�M��o"vau�G]߰b���U��f��Iuu-��(Cz��w��3��U�t��`�tX	Pw��w�ۻ����u�pY'�?��O����״���7���`�R/"2��+��<p">�P^뿩��� �D�ر�-�FS���Ķ�ii/~~@j��u�/nIgC��tW�m���O�~k[qM��p��|��Sl)�T������6��âhwm����v�SC��ǽŒ�ƌ��~��4{;gB����t����Pm�r/��p��qь4+��)"��}�:oV���k�կ�5d����������D�6?%E�U���ó��
2���65�Hᡈ���[~}��(ē- �<�����Z��KP�_��}�{}���i5������f �z�u�_3���jD`�j�����Wm�%�
�cK�*�B�T{����3�������{o��_�/�kԷ�m��~�by@rj dX���9f��?V���)�j<����U�W���yGn}�"n��)p߷���)LcIvx(�<z�{n7A�!��R������I:3�CZ�;Se������.\9J��*���D�՛�V��D,T��۾����Y��s>U�����-��.��g�T7cm������K�nl�8������7s�����
������؞I��ks��2�܋T���v U��!��z8W?t�i��	]m���A�����c�����k�Z �T�ۑ�3�xċ������A��5�8{�?qI���Q�G�S��b6]�7=GFG%ʅRE4�u�J��(�~�|i��SV�=e��z�'��O��xg�kuc�`����-� �=yB�7���i�m�����>\��Mj�0�[�|U	��g��/�0�4�0� $�����\m
r@1�{�S>�d��p)Q��ţKo�������DֱX�i��)a�zcy�K]z����T�j4�X��g�bYDB�V�j[�>��8���M�+�XY��E�)���pM�B�����=0�K��������D���թ%�X-�+����y
�vl����yzH��fl�w.�B�2,����yy��W�/�;._��=���D<[ȧ� IV##c�zUG��LiŹ�]�"Va�G�����j��I��``ȿ�(����˕S��Հl�5���s4^:C�1j-=j�xX���l`�î�J�]9�����u��C��Ps���G�l�҄��Y{��F��!kY�(Ih�fV/�sW#K��GF�'Y�
�n�sV�)���3�5��$��'eP�ݙ�&�lɌ0�Xg�*�Vh׫p��ᅁ�����?g��6ط����]�?�>����,�7���C�+W��n2��3վ�zs{��eW�V�˯>W�f�J���ml+�>����u�[���k��~i$uD_
�0�*G�v�؈����I�S��Z���5����6YLQ�ɀ�_5��m���T +��0_L�#� ��G���K�?�2��w�̈́mZ?��{<��כ�ı���dB�q>�m!M
����~oF���	!		7u���S�e������h$@ ����)1�2e���7����K���ћ��B.�6\R���w�6�#���=:3�h�vcf0Ÿ�7s�,(�_^��q�������*J�T�V��TV=��?zw�GkV���t�t�Иp ����8�F5���t^۱�CAӍ��ή0��̼��L�	����٢�X���A\�f�k��T��\�}T�L7ny���|��Er�\�����1����%���ӎ�ӎ~#���&�W�ʯh��F������6�9�L���Q[�)��&n*ɽtQ]D����9j!_!o��ܟ�6L��X: �3�y�c���-m2]M�Usù�
-��=�*�a������즳@��Ѿ&v���172��m���qc>���q��f��چ��=ƚϩ��/��M^d��z4f7��Rq71Q�Sn�~zӣ�~����N�]U︤�I4��q"�ǿ3�$���rn.M)��}N��.v��8� sI�<#�l�#�j���u�"l��/Đ�R1��c4&Ua��WE���cO��t�qy��Ԃi�߷e��*.VY8N��e�h��%\Zr���mV-���!$�?1)|�zg$��p4�5P�I)Q[�$5m��4@�V��B�CD�urjl�>H�U-޴��?�y���40"�-�V�s5Ux���a�������Z��\�5Z���d_���obݓ(�B<o�D@H��ϳ���ôC:����
a#��T3Mn���V�
�ٱ�m'.�M+����B��/��b��_qN�f'��ݿ�e���j���iޞs�[�_��X�hG"���*N�
9'Z3�B���@6���L�stĕ|+��JD�����U����6� �d����eO* "�����PO�q���L�b	��/r\�	��K��|�B!�������!-7��d�{�t.�`/�=262qto�|�=�]0}<�ߗ�M����4����;�}ů�fx��������%�Q^�^��^�%�՟�^�:w_��_�]ڮ��s掦�ᙳ�,*}x�[�M~6�\XY���D6�2����+2��3��U$1o�7o͐.cy'���(�f��@�HH�ꑏ#���ӿ��B��մi"�1��~��z�����7��t�*�7�#��)"��M ]��?�,��a�,�%sR�����`��k|_����n�6�<[���|��{H�7���a4ͳ��v��r����|J.��[]T(T�v7���a�D�4n��\�nZ�3��N��T&�זS�T�� c�i/�E�N3�svY��PL�"��_�}�a���I+�,u�?���|��f��tVj~U����̒�e�E��=D3�f�/�"w�q$4S<��BϷ��+0yώO�S����c��w75��J�[�1��?rnl_�I4��J(|��|�����i&S-7p4�}�E�ĥ���������B��.�h�!��{��A��B�Ǐ��g�[O�i�I�vA�\/UC��ZH�4<<9_��F��Ī�nH$�^n�%^��"$6�$��K<M&ܝ��rwޓvv��I�c�l�xn�)&9�:a�RҞpH׷���?Y��,}9����s~q���/be�����~�(�Hv�߲܀�Bڐ/���	��艛:�Р� ��gV%L��Ȅ}�c��ؒII9tm�PL� 9C6W?R�g�e��/d���~yl:TN/쾂fp�k��%�=��9����NbU�2��
��
�K�H�$��=	eb���H����%�;W'�����XޞB�)��+��z��j���P���G:�k���� ����K�z`�z��������rs=X�-8�O�@����K��G�)�AB�;���$�0O��|��F�ue����ب[�5�ha��MS;��<�e�=� �P���?�q�$t?"� ���t%�	w�a���M���U�{ף���AЋ�)x߁(o`��B���o'V�8nI�)|����V�-��Ð ��{��6]u�=�
�KN�A�џ"5s��	�F�;l�#��%eY��;��~ 1=d3�C|6|	����� 3����uC���7����Z�-V�|��vy��Zo]��I�r?ؔ3�WM��z��v>~����P��ZD�J�QnsQ��7�<,���Uյ���~��mf�\���;����ڎ���%�XKT�w�e�-��s��p�����`SJ4�5�P��rϦ��i�@>�.)(
0� �*܄������Φ�Z�h����/0ଲsM�xE���A�S(0f&V�fqm5���x=Dti�x�j�W���d!��䑱�	+�7�5���A�������?�9�wy�M�l��*"��vWw�~U����s�|�z��;k��k�k��������?����(���@g���ب]�4�䐇���l�*<��M�"����C���ޑ2�>^�K���~޴��^ʶl��"�% q8��[��>~�:O�0�KI.$�P'���_!��o���˯`��Ȩ����38l��L����`N�����2,�jW]����]5s�������4*_V35��vX~ �R[����B��T^�=�� �( ��Kѡ�(ezoD��h6��R���w�j-Eh|��G�1	�sߠ�t춱Ix��Ro;�ȟIǠ۰H����Ɖ�T9�c�kн���g�)����
�$]͒�<^E<Zzq�w6�����BUTH �ܱW`�8��8�,
��g>� ��=b5%�|*m5�}/7J��R���_��1.��1�k?������"&f�DNcH�����u�+���X!O �v�X���d��r�9��;6��%ڋ�	�Z'��li�¹2*5�)��1D�@V£s�+p�����/8&��	⸒�&�������S!�F�z1
$w�| V�,�"�UEd#y�y��Xy��ӃQ�;�^d���'sL_y�UM�n��$�3�;�a`����Gn�Cs��\�>���B�Q�H��H�=/C<�a%�Z�'{���r�䏒}㢧���-���`����pg۴��
YEv�g ��>]��neS�d:)$i8�E�;��x�s�s�s�d� զ�$���m�`X��G�T�&w�B|�o~휯D�����P��E~dSML�|��}����kW��r� [:~J:T�+�c*����	�k��/��A~���5z��/ʴZ�,[�^��n9=��Lb��VQQGG��J�+JP�z��������i����P��RŇ9�}�����9[��q;��Eh)Ylt2�Q�r�mb����I@�����T$�Gj���륄{��9=��$���DN]�˾!˪5�߶^�עƭ��G^'��"~=��kY � z�$vFd!�����*�߸��;.i������	�s��:�=b��v}������O�+
�m�߲���p^n�Yy��~�L�i�tN��e��`Yj?�0$ºʦTQO�Y�3&\�D�$ �1��zD�l<�A��?�C�U�v��,�e|������}�Yu�I�:�>m?�HR����G�ֻտ�&��2L<J�ts`ഥJX��:�F�I��;Ϧ!5��۔>fJk��7
�.�f��&�/����`���)w�!+���﷙�r@��P6]��O<�"��-�6Ù�K��f{��*A�Ir���,�WVS��8Jl�I�o�ͪ$�p%��b�E��Ap��^dJY����֓1'4��0��;b?W�zj�r�ν(����Ox���M��#q,�}�>��֊xU�V���c5ʶ-�r�?�H8���8N�©��f;j�=�>tܭ�]d���+�5���(�{�؏(xblSf�-nR��Ox�⨧���+!Yg��,s��[9~ƭn�	�k�)G^w��K��a���)�g�{�����An��k[GM��&�/����)	��]ł'�{'2_d*"� �X�3�x�$ ^�����yU�9B^�[�����b�R�Q�D���ՙ���}��c̖��9�/�7o�uOV,��7�t����0p�~2�+�|�>N�:��<"}" D�Tԉ�t/>���cXv��Ę��	�w';��K#h�D�3H���@�l�<�9d�LGL�-��A�Zī�p���i�6L4k���-.G(��턋��^��XO�d��ީg��0��H��C�2��JY��d9ȡX
2I�̫Bb.��[����H,S���C�F�z��+=$B=�e�ɴ@7���X.��ߤ=���b�R}����+���g!tG�0��7ڪQl1��d���wÁߝ�V�5�m�JӋ�qp1�9s��L���A �H�b�%�0ޏj+�#0�a3���-�kC����3鿱�N]7,9��
�> ��&�/5���&52��y}0{ee��#��Hg[��ͣ���#���B5K��(k ԋ�FC��h1��ԶɄ�����_��l��y��Xq^�б(�߿�����P�mRc�-o~��ZX^5��=6��5?�hm�>��r��qd�F��5��û�b���û�F���0\��1H�����PY�H?^���Cvv��c]s���.A�ђc�eI?�{钑��cmm3}B���򢍟�:	�"n_r�v�(I������Z�@�ud0�ʟ�2ea������Ȅ>�X�ޚn�>?�_MF8::k�����b�D�b�|F�c`���?��-�I��q����j���|	���,�T��׉��ꬠ ��SÇh2#��x�h�/�t���SPe���0N}��r?����cVb<d]n`yY����Zj$�R�'�ZX?a�Pja|!�i�a��N.��u9�C�5.v���<Y/�`҇�j�p�gp�E~�N5ӥ䌩��T����s���US�i�ta������ݽ	%�L����GY�p�be���78,s��@�ӮO'�����rI��9���;2���S�J���w����V_��`,���'B,HW�>7Y����Ǜ_\s;�K�m2�e�a!�5�M�Oq^?v�'�ݜ^�~�|lO%�raQ�K\��=>�ւ�p�*{J7���<8���ց���2DeS<���o�ۻ$^#;��;7R�$2�Q�I�!���c $��9�8��,���� �r�b� nj̉W��O���+�9�{Б`U}m-�t�ȍ��Y��������C��z?���O�u��y�?�p�{PBܞ����ԉ��N���#��\�+��a�(�k������/���Vת��|���̹��v�G\�l�r����`,���V�L��q��Vɼ� ��U�	M���i�3i��Q����`S�a�s&�}��U��9����I�?��˛'+~�W�	����skG�a!���I,N�v��	�����>�9�%�BG~��$�e��^GA�������6vG�+�b=&�ܩU,��.4��|���),��ia����E� (4}��PO�6;�	'4e�L�喤���OA�r"�M���^�����
�AȒ������c#�h�;kJ�k�^�vE�,�v7�4צW�E�lS���=N4m��$,���4���rOO|��?JL���ɂ�C�nO=�n�(�}C�4_=�����Q�S�ZL�}����>p-���?v�"w����7¾y��Q?'����5?k^���n������0̀����M��OƁ[f�tHY��o�*�.��X:׃�!�P�
f	~gbf���W�d�^`�ϯ1@�:�-���#-;��� Z�� �q��'&�������u�_���vK�D�U����~�q+�ߧ����,y�̔�w��g2��O����S�OV[���k�=�K��GM'�^;^z'�^;�^'�~�aK�����9���-_b���C;֫��ǃ�*���03&�q��.�,�H���(��P��x9�.��S���p��04�r���g�����*k���x�?'�WZ*qk�j���P;�Dq��mI�������e)fFeB뮥�,����M0;�{�X`Z� �-r�����O�]�|�S>�%���*������E>��Xq�S��v�5v��������U�`=3m|aQ@�q�=����\޽�e�|��+Vމ<c�H�3��h#��ZB��#?ܫ!��X�J���s�K&L��^Gk��axƮ.N̬l�y(m��T�	i:�:��W5��fe��2^���tTm��q�fw���DTAhm����MjǪ'�Y��ZLT�j�Wo�V��5�h����ߺ N3ȴC&#qz{����v
�;����@=7�\,��ָ�.�Y�##!b��%��FoET����9�~�=����a�^-�9	�0ڰ����,�p4���X���F�.��l|E�?�2��8�fq��}{�'XJ-O{wi��;���n7�$~���Mv�M}��1�_(�\V6��%�^V��@S���)���6��s쳰�Zx�I�E5֨��;}����D/ c��>��I�hi�V�ʹ���f���T��H�GDj&�,Ca��b]5��j���[�e�uϤ>�L��U��1:�mPhZ*��hAc�1��[a���3�����������U��ENsluY4��}�����iP��Y@\`�Î�並�E�V�V2eE\�"�a�}���$�,����,�vG�z2��<��k΋:_���vw���?rt^��u^���e��U*�o~���Etp(3�Sʲ���m�����&I܅H�_r���� �D����R�v��C�V}C��6��O����e�`�ilqn: n������5CK�� zi��}� 8����\ژ�����PEJ�R��=�P�~���f��i�PǮ���%J����e�����E�G8Ӆvj7����� �#q��^�~�k�t��z*�7MD|�Qѧ��g⠻��OA�A��b4B��ya�0��/�w���3��m_����?i�K����t���x������ؐ��ɗ�ٞ�y�"�2*u�5�A�[����5����ƟE�[4����"!�d�H��q+�h�k#)̂��;m�p�Z���6�<�8��/<��?�z��Ȳ�EH��� ~��a�7�>M��;�c���'|Dz$����iP��酋|�E���Sv�j��x�������~�u7�<�p#�Z��vx�������ӖnnI�-+�T�iY�<���xg�n��"^>'�{X���[�Z�v�K���;?U�Wd߽�]�������+�Š%�ê�o�W��A���04ɰ_l���¿�v�q�o���r���|�k{}yl�Yt�z�H%n�RW&��9��c����v�W����+��J��5~q����o���eNc#n�x���Z��h��y�f���k��	��e����$w��Y �{X>����\d��{)z�s�zum}���lV�Q��
v��P�S�����?��v�����`g�5���q�S��ٰ���:�7����0�sz�\C��>���(+�	�҇����ze�^Q�LR����~&O��E�/�L8�|��*zy"�_6k/�cR�^��v�~4�+��|ta
���lc��x.�ʢrI�t�[���RAg�ɹ^���w���n���~1ݻ�@Cֱ!�9������d���YպÝ���6~�1����y����)NE��Ռ�d"C�� ��
Lؚ��l�٤%��-D�a��G��l�:��u��������O2(��q�-G�)���b,�%ڴ�i͍'�`�R�@��'�%���O��M_Դ��ի�^�>P��N(�ss�ƁL����[<��QVͯE^���2�{��7��U3W`����o����nۼ��ɪ>�=��tœw$ѼT���@<��ʥ�;�םγ�����_nZJN�+ׅN��y�B]�CEeemK�Ҕ
w�~����d����
�Vb��آKʢ-��c���g��*��,	�N�8���s���Ȃ���<z{|�������/���P��}jO�4J�������4�u�6L�Ic! U�1-Y�d]o�M:)�ѓ����(���v��3Z��`��[g3��\@����J!r�+ �2q��cR����~�'�}��34Z|��*���KpA��ޥL(a�[������֬'�9�:�lB9�$n"'W}�y�T~\�jVj�c|j���Œ�����	��s�"�.M6��k`��>p�p"*⧷�w�t��զ�A3�8�tNw7M�R[����AZ�^^ޑ�.QAƄ�݌�Ls���+ߑѱZ�M�K4�����7�26&p��bӕ��,�a���z�>\^�C8^����Ø�y0u<�-*�ӽI�\��e�L6�u��>�NF�ڿfg6��qL_+N᝚{yE��Rh&������������3�lwl\�� ��6�����rp���������(���k_n
G����X����������60XE����R������fR�7h�%403�0�Y�{�\�<���\g���~�N&�o4�soO���h�myS���	3�J��E�J��3����'I�+Z�3�4c�x�+�F8��e(�?`��}k���6W�;�Fy�|2�T�;��7Z�t_x�s�Z+/��]2?W�ʯV��&�˳�22<-��u�FhBi_�������TI���FgО�����-!�G��5�'L�	7rqO"�]c��pʙ�]߾q��:�mQ�h�#���r̜������|�h��ll[ۻ�m�֯��1�dc�Vc�v��n�/��}�}^���s��{���	�t�����O��#"YgS��������2'�,�b�7��	T���\���.�U�eIR��#���8ɐm��.(k �����Zw�g��j�����P��l�ٓ���MA�&���"Q��5����N+�?�VC�ǘk�15s���Q%
E!(Nh�$�b�i5���L�C���,�}�pm<bM�s���M)�9Y ��b�l�Y�N������j9�d�W2P�t0��e
�p5�Z_2)�4�G	ڻ?�XF'?�ZA�f�|N�2zm�hnQCl��%�S� ���uv���uē߈��͂���QvG�Ex1��5&,�V�d3J�_���RűK�gv�B���(���T��fq7(���؋\��*u[D˖��~��P�/n�q��ɱԈS$Ƨ�'��*�30(�E���n~�bR�����*������*�	�S���n|^��>��T�G� q�!�LIj
'��Ɍ�u��<�{����F����|i	��z����<��� t��-ؿ*n�è�@:1/w�h����FL��>@�|�so�?O*�N��\v������ɜ���Xf�	+I��g��Mrm���ȓ���Wo�n|��vi�c/�T��ïL/++/����~l�^�	ܙ��A!���3��V��+��beQ�Ro�M��{m����3��M:��3Ĭ�	���p]�2�-�Hj%�h��,�Ǚ�f#e�q<c�I��v�L�lZ�ˍ���).~�nM��YFAO���a"�Br�Ybt�f:�Cƪ1�~e[�C���e�~i�l�j��ުi�cUN;��5�'o:��������͈hț�������=�W��XF�*ڱ^(N�?~+j��E!�1I\�Us���?�O�
�h1��Ms���@A��J�@̝�cim�;l�G���τ�n�3�V�NGQ1u-$$�tFF�Y���PY):���v6�i�e#�l�j��mmS�h ,*��K5F�����g��C���u��?$9���x_Ơ�`�&��f�*[}���j�g�A��;��fS ��Bq������s6�[�]������W�)96�1Q�\��8d6Tm�������۫��cwh��}��f8��f��<s��~���u�U��|�|�vD���E̴��"9��=�+
���g����3��<��t�non��.�d�L�g��o茶b[���ȗ�<Kv
�8$�W���t���Ω_�J�۠'�;onT&��j��j;	�#��G���p�h�J�1���PK�%���V��D��d�ͦ��G:�T�F���3x\T;N�G`���w^��>��������@�@OFFF!���5��5�����`�];%t�c�� &Z���WI5�̣��P�V_�sG�si�H����h������F_��I�W��Ftpp����=f����-�o�S3oNOO9"��S���^y�g�OXWӍ���˨֖`��cnU�AC���*梺���TF��L�o���Q���nb���m=-#.�Y>T�����iY+�����<g���-������>b�$��GF��UF�����`9�219�*$4����q�ŧb0��ӱp~��!Ӓʣ}��(N����<�ilh��Q�$#��_<Ӓ�uX�#oק}�������I��B�4UY,)���4�w~Σ����������_dl��"�i2aK'�`-����Li#�V�bY�]O�?L�\��j|�ᘖ�z����X��9rdXD$$���f�4&�lܲx�|��Gf������H���)^�C�ŵ����v_	�1�
&t�1���H���2�!�F�q
0|�<�5O����� (��Y��%�{l��sA��M�	��ˆ�EMMZk�*.F�9�Y�C>r.en\8U�/����{����'����t���r�c�,.���M�w��i�g����L�88��5fÔ�t#���(��p�hL�1v�C�CZ�c�7�����8<��*�!��9�ڙ�ց�#:]���b���B�F�Ѵ���$�&��{��K+Tv�=�&��fƐ���N�Xq��P����U5E
��.�r?��2�����Ц"��0�3�J��)Q�
�Vf-�n�����a����k�+��������S��܍�<G���(���c�B�=��>�l�;����C��.���ۢ���}:�J�|�� ۩y���	�����0c!�~�6QϪ�i���@��g]�H)^���U([6��Ϭ�����lL�H��Z���Xjux�t�K��R�G��	Za˔]Z?�k���'  �[����´Q57�QT�Mp��Z�u����@D���U�YK|aiF�l�q��3YBK[1��w��}rr�#�,cpE`4��>��X���/:Y,�M�}�%��;>3Le�I�����7��� ���sV��ګ��ў��W�'���!����L�#e߼�/+T��`�˯/�H����<��f���X���dcU&�h�/���(���}���V����$72$%�H����L�"�vf�1��N�[��D���Ջ�����w��I���w�� K�hr��oTh����h#M���y��l�H#���S��
{/��uLvS!��O�FN��}�7D@�z��$�Z`4�p@�1E�8���� -S����U��ᒪZ��
��`�u��i��)d�.��yE?d�^�J6(ny�)��x�յ��~�f�W�,�7�,_gPƙ^=�u�Y��,=y!M�ip�	��������n?u����'G�i�n�֦Hx}�^=���+�ȗ�am�R�}럞�m�}b;��j�Co^Dk�!$,�	وQY��d�@_�Z�pi�lU���4c�����Qu��(5�i�YQ�}��ߪv!��M�u����sCf@�\CA#�Zp�}�O>��k5�KNl5n�}�2B��R�p�+Uo�>�ZaMM�IO��s�%w���<YL]&� �7{�x������v�3�%49� 3�<6{�n��z˫�r�N:� \���_>�.�[����P�T/�<�~���o����c۲-`�H�,��
ι�&O����A?�ϕ�H>Kp�	�����&Y��Eh���p�>žH�i�p�lʮɪ���U���=��H�h>g��˹}��u}��U�U�ne�ś] c�F���AW%�ѱ�I��^��DXW]�'�ݢ��	g"�pL�fb��o}k��\Ka�<�h�k�L�֖�ۊk���ȉ����. �p���LQ}�71Y�R�1�!�8b�ǡ��e���?����f�n>3V��nN\�ޯܮ�<���W�����N���j���a�U���K�zw���v��VR^�c?_/�AY��شGFc�2���1O�ʊ���IN~�5����NR\����A�L-��y`��]���4��H?|����r)�k�x$����bQEs+�������O'�4�ҙ0!s��4�P��<���83|&|P�d �@�鋼�n%�RwDi{}	�}���lQ���)KRjV�aAY�������-5�� = �v�f���V+	�.곒M6�E�&_��#�t�FT���?���kh�x\|�a�3u��s=m��Ж�]�R��@�z��@�tv�z;�z���xZ7��Nܻg�t׃��b�ElԖ���:d$��W}��b`jM���u��W��+�Ȃ{�z����u�ʀ�R�{�6�6U3ȟڊ��?qu����:wl9��EZ�)�-��	da���űn��*n���j;�/�[uk'6xڰ��~ӻW���`8���O4Q{��PC�x�!�Б�C.�oG��*E@�������jnO�����%���mަ'K��ܽ�49�h��c����M��	�T̘�Δo��Aר�?�)��mw�S�Q��X��}Z��v�*;d2�3d��񚞞uk"�Vi��V��6��"qߙ2��/<�he���u���.�1�Xs���"4����1f	��:��+8;�̩e0⹩��;���N��V���}�d ���X�ZF�Q��|�e]Ŕ^�X�l��ߥ��`�,8l�4�X=��%��M�LY]��4�F�]ܽR1dd�Ә��Ì!7�7h�BmbԚH�����������N5����a%U�"���c�s]���ґ�q׸��wm�;H�m���+R�q}��L��P�Q�X�#׺�]g��H���ЍKJR� D�R�M�d�&���#�&��VO�h�QxRe�S��CF���E�^�q���PE��]�:��y����=j��(e�┑�`я��ˊ\$�a&�iA�X	�L�A����8���P2��&
��k�M��y�sq���qS���,ۆ/�M�7Z5Ru3.�Eʷ�5QA[Q���[Ӵa�Eo�E�W�y�䅢.o,��~�����|mX,)�P�h6{��d��l�ׇ���W�b������KT��s7|�!��<:N���M.�p$)�6o����&�)�) dh_�d 6Pl;u�<<^Z�\_��w���
�l��"��z���kM�?_��2�F�l�li��y�E��\����-GMq���J+46C=�22\n�l�����*�ے?��?e�/X�hX�çln�qj���(�d���A\$د�:0}�jj�}��$�J����Z�H�?���%@)3_:=�S�^"���lF��U�b5U���NW�[}�'�,!zF��IPf_|�$G[k;�it���C��q�g�	��������V{�oE����"��sܖ���A�����'> 3!Bĕ��-�o'�'8�P�XP@�6N�T�>'�M��|=��,S����N�)e��X����}BW
���� g$bn�Y�:�j��a��S�[-<o*�
�)[�L�{�aM�F�NA�y�ѵ�e�GD-�G�¿*��T������Vn�k:5��"�a���]Ƿ��
�~�u�SVV�Cz�jU�C�0��M�-P����}�c�]�}H�)t&��2������?w�(�Cۿ^�L�_�/�̮*{Z���^2Z�!���R���*�Ȅ���;ë� �*~%SK|�V׸�t��	���w�S|�r��dʃ�
KQ�p
<�u�G"fx�����6G�	�)]^
e��������܉<�vSd>��a��BRN�T��l\=ɡ�+i��ضj���0���� iga S4��D��w� �RI�7��A/��J����,v�f�*Вɚ��U���E
��v�t��#��v����v��4�=��I<%5�d��\�8��:T�2cl��m�vC"��M]���[̽��n4��4C� � �ŃTہ�
s愈ߟ<��j��8��ǔ��3�-q.Q`��(��$M�7ڇ__��]�Z�kȉ�LrT�O��
{���������W��.ȉ3�~�P$j|�,-	R-VҮ��F� �М"��$�B�l��dg%�#�]�~E� �(�emM�J�>vî�{%||6��(�E�qs�:���3gb֖C��7������r,N�����.m|���g���:d����u�Q�ao�eF�BRU�
��3_�ZQ�Ihs,�D�KLJW�b��jP$�rav����&�$R٥�%��Ǆ<+̂W9CM��7I��Xl5-y�m]��b[aW�ׅ��Y:��WP��p�LCG�k�OC����u,zZ��S��4�a���5Շ$�H+���s����ʮx�������r[	~�	�ڋ�%# �c�l��^#n`� ��c����m�:W(�|�aM���`��#Ie</�*��kc��Զ���+��E
�*���0&�˱c�������E	��*W�5E"?���?V?p�#��Q��Q-Mn�xjHT��@t|� ���`6�޿�*�qj��c�*E�� �u���|�_z��c`�v������u���DF�|r�Q���;J��?m@e.�(.H]������'�]L��s��P7���)��Ь��1֩S�`���H�Y1��<;����O�(�U�r~a�4��r�V��N
��|Q��3�恪��]U��gnz9���n�%��:���������(s��1���9�4A8i���-Zp��i���BN A-v�XSD�g#H=�C���[\nmu�pw��>s��:�<d�Q�I�����M��O�_�Dq�JC-��� Q�WC�3y&�MZ;8�̖�����y.6-LL�=��e���F�T�˯��2m�쯞p�n�&�vc��-�;�۟��ȗ������M�95�sK^�
�E<�
��R���_.��ƋG"���>���|ڲ ��_%��$�r�bI������R�>��� 3O�z��BO{��sb�����zp�aT�f�&n���h���.z 9&5g��w�7�D���2l�E�`��7G����%��Ř��ƞ���4�K���D#��[��k��I�
ל�-Fe�^ޥƢ���Ί�X��8��P�S�V���L���E`S�L�<�}Q�!ġ^\�T������ݱQ:Q}�h���	��J�N��n��߼����l�oi+���馬p^��Q����K%�}�O�z�iY _�3R�8��|T� 4gȚ��N񾃻���Y�`bI�i�c�%�iʔ�d&AŚdh_�8t�+�U��XР�9m�-.E0�H�S5�8GI�׉b�d�-�\��)H��zMZ�⯑�[�{�E:.�FC�PJs&�A��Ҥ�R��1M?����P�ն/�x��7|l���N�p���U��rO> z"�or'\"�6��1�#]�F�ˇ���yIܮ��V��'E:��C{����'�y�����izɏ_W�D�E~'�CnP�}�U�Bw:���T�����H=mР�������שG������Ih��ְ��3;�5���;v��rI	�����S�����[;b~y���N�7ᚲg0��\����$c�+���'������c�c3�M_��#��d_z�Q�ߟ���/��WVWw�fi|/�C�}c�æ�j�^l����1���{�b</��Pυv���|��i��	�'(T:=l�565�͂f�\�AE;c���2�1�(�F��aN��kj��E�d�����b��.��כ�aI������d����>,�/�!�G�������3�`�p����;�dШ��w+n��`aC'_�-�W�d�*����*�h&��`�X�QlN�Е9G|�)f�'�K	�J���M����ΉJ�%�Ȧ��B0#�{��9�i.ӣ��iY��|��|�a#���<%�T����J���蹑#>� `�tG�WjB�|�@o0"��,J3Z
#ъ *�P����f�bu�ۿh	��X�K@�ZJ##��78��W�xR_�yg%eΚ�i�i/�u�����i˫�-�m�Tj�}��X�>�2������K@�Ն��I`�b8��2�9H�JOR&<����������mw	�gm���l��ѝ��[f��Ғ!nl5�r}������O��T�"�r��?7y���?OKQ�O3ћ��I5�`��	�I`�zN\�g.�*>
�h��.�X6=u�x��1C7��/p@eފ�jQ����ԓ[�G��`ZI�<�qrQ���n�M�X��NG��>N)"����Q'P59pR���ꫪ/�D��0$$�>��� �c���3���2:�HL3��{)o���=Z/R5K�C����"�6}�t��(�	C��2�We�Hĕ�8�~���A����J����z���d���;��^-cB��Pخ�5t�|���-�����fi�!۰��%����J�MyUU�aBɯYj�P��A��i�����l��-��|�"c`x���'''�I�TYZ��<�v=ڢC�f�ٗ�@h���s�¹31ɤ�V7Mll���2�x�2��w�wm˫�/�d��f�� rb���u�;�~������?��~�G� D&��x0Vv�*�w�$�D��s�f��,9�9����P�� Jx��/��U���iyc���#�l]�핈����⬶a���!�b]p5P����݋-	^[��O�gJG$߫ _�^c��Y�����2�V�Y�O�:���[�卣��M#�	;�Њ���S����۳��Bb ��/R�4Y�똎G��ɘ���p�2����1g�j�)�I37�5ԅ8���� �xm�h�[� �#�����1h4}�1��G^���]��y���ȢxZ�<`�����)YB[��X5������Ս'�(Ѝ�3z-����=�����eQA���(1�0�emH�������8��9�)ĕF7pu*iԉf݆,�nnI%~�p�?����]v���v��"���W��x�*����h'MBE�����r�ɁH�l{�Ao�''6o��|�D.�`���a�3���6�#Ё����VҼF9��I�+Z�Ї�L���Y�@XьԨP���iQ��Q��Ual���N��UZ����G��qgo���`�;4�YJB���*��$b0�7T�?�D�45H20u�1�	�|�C{{Km�VY[�7"7{��IS�`w�A���f����L)�!vpq��AxK����/>����c�
aS�B�7
�:F��^V�L����6wPR���}�Z��!���-����W�Fw�U]��#�!#;�����f��%E l��Bhh:/�@53p�(>�X�g�Cx���$ HU�j�P��Ϸt���g�l�1%��g2!ߩ��Q��8�����O�"���Yk�'�j���W	B�Z�z�6�<2Y��LR��
��P�*����e�m������֑�"��%C���3������U[[�ښ��{���U�S�:��������wO�g}�.�M�K�tP�a���'�>;gc��Z�M����.�S{����:�B���}�|�؂�����o>���� 5� z��'G~��@��1�i�IK��{"+�ǿ�����T��Hg��	24Z�n�-ˆp��bLb�V������S��mt���h���ǋ���wM��sƐf�ʀ;<P0�xϰq���z
9j	9��l�9��?Tk�+X�9���~)*��:��d0������gmuF����\��_�2p[�����pC~W�U���GaD�#���ߓ���Sp��
Tp#�E����������X��f�]A���!)���Mri�9o��˦qU��U������,H��D����h	��P�ZD]3�֛��$TT0�k,~}e�7��ް�!2��6����u���+���Y�2�h�y�#V�2��[F����|�A�E@�E�ŋ�{�f��"P	��vȈ4�N����T ��C`A}���F�����@�޷�ww���1w(g�	��x�%eU�|]�>~�*3J�#���եPV�ݰ�����~~�M7ۡ$��YN7r���fdg����Z��Ǆ���n��؈r��d�ՖU�ڢ��AS��b����]W�`���BF�iym�x��k&���� ��-�
�}v�!������)���Mޑ]��)��,J��߰T[P�nԴ�aT�\)Q�c��M�<�.{Q[�OlNd#�o�MS�H������]�o��E�,cg��GX�D����������C�|��ف�#���c0.��5�LQbn����%y:RQxV츧K�����fˑ�86~�0��4�R 
J�f��ӷZ���LI�t>�2��͡
���Z<8_o[{܁	�J	������Q��9�^FF�������CQr�!5T	_%z�N���V-M,�FkR��j�C�;vp#��.�vo8o����W7�J���ˊ'�m�L-c����� �G�,�)�����������;>0�w|��҂�w�X��y��Y�Ȱ��4dˌ͇����t����� ��DpE�C�����(�OZ2n<  �?x����C]u�=��C�W=j�xJ�?���Ԇ*���؋B�`T���찫��0��\�f��EU�����+z@��b�<�$246���[�LZ&Yᤛ>zr9�3�M���4�A�;�{�$�	f���SZ�������_'=}���?��:��@Ԁ��t.M��v:�,x�)Q"8����9{�Fe�g����_�x?"�U��l:�7��B�"�a���z۠��~�ˢ����)�����gG8(�����I�N@��!�O?��������Px����L¦$p0,�(̆,=�_�}Eؠ��K�-��>��ȁ�F�������ߌ���d����}ۯ��4t+[]E���/�L���x;q�\l�p��Ljwb���V9�=���`E�D|��+���:�~��A�TS���g��+^���L)�>�Юa6;��^Nq���0o~��pG����<-@bI�~ƚSKSw/IC���cz�D���E#��`���zO�_5`��H	�}����rov�@���,DawiÔ���h$����k��Lw�#N��D.����Ӂ�NG�TU�-�6�c�a�4� Lg߇��k0&��#�8��-,.�	����,Mi�ާwh���Ns3�D��c�������P��(�GV�KH[��B�-<��>����Wر��X޹#�n����ˣց����c�K�'���'�l��$�6d@/M�����,<O�}��x)��k5�_Ml7�UC�R��ע<�@�U%j�]�5.0+�''�� Pf�$�8���_>�Ǽ?����}���o;�yU�:�fBjKF�Hk�mnE,>e����M�ߣqٯ��'�ZJ�s8�Y�K�S� y)9^�@ox=�m�����j]����P�+����^J����BO	B�1oc�?�b��8��Q�o�x�����9y�
Z��kX,���7���9to�%I�s��!^�^��k�W\�����y��f+=d�'���;��#A�����+<�۵r;�ȥy�B ����v���]>m�<�0:B(v�a#�M�t1O}�l��tᮼ�5IŰ�6�L|K�� �ʹ �7��� �@�--���0��-��59��(s`t^�>��6w,V�t,@�p�d�>P[�n�����C�3}
���i�Y-m�QDi�$zm�A펪hI�*�6���取6��ʛ�P�ڶ61V:Ÿnuh@|M}���C�]W�*�� Vb��x�V޾�*��*���*ݎ�j�9-�a���<	ۛc��N8O�l� ��T�V��y���M�Q�M�!'����.Q'�?����f��Ba&��"n&2�^"f}���	u�=�6_�7���0Уҷtu�,v�)�w�>~�n���y����6%����N�F;:4Q�IL�����vA� '0���j�t�K\��*��݇��a��麢x�{� ���)��'�JDh��0����$T��߯;�z�zS�}�E<ЦF8�	A��?��Q��gd�p����7��bM����o����%.?��g3���a=\l~���|Ttj렂�����sX
�=�L�'�����%� į�D�L�$qR
͂5p��CO�a�Y��*^@��R0h�k�a~�s����ǹM}AǮP6V�7�:��Q�RՄ���-�n;����o�]N� m� Ƣ�,�R�~��ֈ FC-Q������u�����u#�a@Py�nS�I��MƷ�=w)O�dJ
��fLj�����777�� ǣk��j�\a긼�-���A�ΗE50m{c����3��6�r3 '������}�F�®�*��������fa���B	�g|����~D�,�y��̱�����<m��'>��W�WTD�ܢ��8>]�U��8����S��MF�Ş��]����Y76P(���Uv穎Y�	�9#�cK�c�1L���hkI�6�RJ�ON|��D��p��#L~�.|½�&��A��|�K���Z�E-Sp��^�;)��~�Ff0_!8�Dqc���;k{mً��Mr�ǳ�	�}#�i����ܦas �"r{&�;�ƫs|v���9 ��颦�F.��,܄c�8�[ѐ�k�8��9��i8��s�d���d�I������گ��W�4���`79�'w�����1F<<
 �m�V���l����=k�m��s�Ѓ*��:�<M��yF����(2�8���Ͷ)�)͠�ƴ�{����K�@��@�	����҈`˯>�T��+mAO�4��"t����+c�F����q�"��R��%�E��\������Tk��\�I�
G����y�a�1�iŇڜ��l�r�
��0L�Ѳ�d��0[�l?`Y���S�I�"-4Ϙf��LF�H����tR������I$��:�Z��%S��M����__��g	BӋJtWס�XJ���@��Dܐƻ�o�.��l��`��k�����f��=p�a !(C��Zx�h��� ;��&'?bx�(�=�`��q��{���x�g�ؐ�}+�Hmlj
�"���+`ר��Y����!�����upR�Y��jdO������w���V�]
���ckk�7���u����X\��G� 9��nh�N�P2����ݳ�=w�a�l�e�O'Xi;�&�)��;�q�7N-�*G�]ر��s�Q�ر����m�������m��QN>,���λ�[XX�yr��F[����m��
�Bv��O����<�8�0}f\/&��o�t���W���Dԛkk�L��~�O��{}DZ1��n���`�	��VW��
�Jߖ̸���GhΡ�;�4�4ʱ���j9\�=-�a��E��Cvd�d�D?u6xk��؈��0j]I�yq���@�����Y�u�S
�TO�dۛ$?��;�.��mD��
�ԗ"Ux�_E�
Ӄ����B!��K�Ù������k����q<���-A�����0�QK��L�e{���~��b4# m�o@���0�ޅ{N��ĞEe�+Ѽ�V�j��h�G�E�9��&ե�j�>���\0k�W^�*��@T��ݙ��7��
��-�+t�ҋ�~Vx���,u�m�0��P�6�Qs&��K��86�v4!B�-�>D>�� ��B�q7(�ҁ����T�&s.7*�Ƴ�΋�a]� ��gii.=�H.�<�g�I!�`����!��O�)۠n9+w��kG�r`�"�Z����'��S_ӧ(ʱ�"�'c�p?�4��߳2�0?��h���
��P	��5��P�N�$;�:
��2h �0q%7���XSB��bM��������ŝD������߿qΔ�k�Ǳ�Ę��[�g�D'
-���2,,=�z��;��=�=m��e��JX�e"=�G�}�݄��	C'����ݞ��G�yytGuAȼ3�L�]A2����4pn}�p�1*���Iq��KH���X������R6p*�D=|B��-�����>D ��M��Ch������T�.I�6�`��9Z��џ�Q��/���nA��ݱ*#�e�� �l�h"m���E��%!�G&7��?�HO34� �1�Ȼ�X̠��F���/�JB�iX��(S	k�`�,�pE
I�A�Z$*Q\~V������TW�{�m}rc��wE��,��lQ_��f���C��!hG�b�jkԬ�D��˴o0%�X���h/,z�[:%�j�a�� ����6���I�>�^I�9�^W��^�;.�q&f����B�zB����/�~S/�
'LS��	����Irb�.��5�-�Wp �(ڊ}��mĆ�I)e!���d��A�M�`�'�� O�_F	��#-��(6��9�!��x�?�J)�A�����S�!˸,�0x�7\���'T�gfT���B�,���)�H��8�M&s��$�0�' �BP� -����6�x�Fr���y��~LA��-��%!��6������s���8u��`������Q�����R��-D�E%	K�����G����KJ�I�P-��h���Z��|>��[����}&^w$;vT�ڶ��?A�sff]<mh-0M5��0��4_+uW.�璾�⠫J�VK5��ecD�Ǎ�����h{��Zm���Ug"BE�J菀1F�l�������ȟ_�L��$��n]�e>�	:
�T�bxK�,��.�˻)�<��-3c٩�aU:�m���J�O���#��-�G;3��l�|=s�	x����z��z�x�z?�zSy�z���s�u5��i������}|[��.���3|d�D������qD^�Vb��X��6hL����o���%�@�p��s���w�W%�7t�axa	��=n�l1��=���{qy��ƒ��0:,�;h��U9��`O�}֒J��z�p�T�J�k����U���k�8%�.��R������b��*Fz���T%诒��ߨ݌]�ߴTm��YO���/V|�.Jtn�ԣ�P��0Sa̞�s5�ݝdx��d�m�%1[Q���s!�k忞�M'RGs]��I�.�D�s����.�rW�S(��O7��ʪ5Aq��NȒ�mlC�L�����7�+�^�>Y@?�®%?	��߳&�.��̇N�O��Y}�ՐwD�q䴗��u��RO���	蠻�ɪEo�(ѽ>�܋y����=@�|nuo{ubd�h]+}�=�ǘ�2�<v/��l$d�*��R 7���G�ɯ��hD3jQ�&R��d_���k~����˛y�.nIR�G<�dmT�a��4j@j�-��c/���������Mǅ������#����*��Y�lsR
�lYU���I��J��v.��7	���t��9����\�b��=���9��0E<,��b3��"3嚾w�Mו�~?_Tf���v�9��R�7��E:I�):�,�t����H(�ȡ\tɬʻ�eLWl���r��(I.��Z���� 2ѷ���8%!�,��}�&��_;��ԲD�e�r?�̉�Ţ�.�sx{&��XDZ��" �iG:/n��M	�Zp�k"����P�]�'��Ic�]J��6�b�(^e��o�M�U��l^�_<(B���L�9H	��hb.��6��-K��*n����-ԉ�c�ü�0�Z.�>���D`�����=�P��ڊ �>����Vmp-~Bx��b�8_x�S�ژ��D뿱��#=i޳��B|�X�B��dÊ/0goǘRL��\���'����[6#.XE4�"r�	v����!.���"�i;�#w�����>������,>��e��;Қ�w��c�Z��л�_�$�bU�i��A�B>ov�n�O?����26�\:��NPp���˔�Iz�vU��L�M�?�I��Z���� �Z`��{8�r>%:D�O�/��k��<���N~*(��7�a4�~������������������ e���&Fm�/���e+�����M��ZƢ����;��a'>��ܝ'�]���Yc$0�y�]e�h�#��?j�z�Z�g8�����؜HN�*IGd�7^�['���_B�H��N���w^�q�0��d��Gi��T���q�$�1�<�y�w��a~=i�;��U�������-����2��& ��b�:��Due���)�u � v�%fxH��axl���՜f� �z{�:.�8�����T�����I�t��)]o���q�ut��NѶ�-�G�YOc-��lw�~_��{���MQc����	�$����"ts�#5��������#Q'�C�0M	~U@ǂ��R]>�
�f�(fn̂��Tys�Z�o���Sf>G�`���������4�F^�_���Z"'�N��P	FE��Qzj�a����82�z4�XO��@>J�]�p.��b�7���������y�-�G�'�0/��A�\���#ZE�\'���S�ؗ?B���)��@bu�/�m�??ы�X�#�����)��&�F���GF<���B��ek	B	��/H��$!���ë-�A�C%�x|8�f�DJ9(�N�*�5����ᒊn(���䓾��Lqozh�W�V�������u엚ի�X'=�NL��7ץ#���A�fA^���:`=zi�����z�ek�h,�4Vi_A���U���l��.=�!�W�aL.�'O���(�a ��K��1l�q�r�²W}��a�E�������/�=ڊ��W�Av�PE]��(e.hBӨ������q�Փ��!A)���o]WS(C�ůtMK�F�����a��]�Y�#�@���Oe%Cm�o|��`��t8Q'5^d�Y];c�x���Փmr&���Dje���^��ZkwE�|�~	}�n�7��[�����W���^���zQ@��-�<|@\��-t���L/_Ɂ5$@mhs,�:��UZd�p��R!�"
�}+~��X�ʠ8��������	n��n�\��,�h�E��Cpww]􃷾���3;==}�9�{��A�A�7�Ҥ>1C�}.J��b朐{ݔ:8:r����!K�B�����fYe��d�Q�{-B�8�5#?U:.:�;�zϢ��V�o�Qܓ �Ff���勘�IR)f�8�B����v�R��P>��2j!@9�\.��1��&}
b1��)�NK9f�]�F�_q����ඣOz^`mj��ݷ��s�,�������N�P��#���7A�x	xxZG
�?Yjbt�cU�-i�yx���F�JN|	g
�Jx��s���:��Ԁ�"���H�ŗ4��*����岚ӡ�u�1x+9�Q���ν�n��C�#��:D� �[럿k�w*�p��,'%�o�RE!Ɨ��x���Xs��M���&:����-�~\�sK���F�Q�!Ioɗ����ΧS�ث��!���e���c t�� ���wO�?<������#kR�x�����@f�ȼbc2��j�~f�#q��Ȳj��
f:A'�j]
���K����g�|��0 �A�J�l��8����z�-��EH�}�
����݁��$�:�d��H�I�@�hJ *��/���������\�Y�Q9�I%T������9�����n�օW����G��.�'��;�+o��c�x'�Gl�����0n�;�&��yTx���	����wv�ќ���)�騒1�Co�b�W)����V+!�ҏ���)i��O%7𺍩�Q��]X;���ó�����b�ZՒ1�7Y��C�/QY��W���>�h�����*��;��+b�wu&��^詐r�qו�me�v�ʆ�Z}��Q6�ǵ�O#G�pd��/�=��Rt��mө����3�?`��^l��n�YeEQ�
7̘y�R�����V?��W�ꃓH`��?��r�'
+o������I$!�S��û�mMme���O4*��_��?.bgh���ռ%�$�Μ���� >�c4C���{o'-Iamv���8�:����:�I��~-ȹh~�K7V��^�y�'�uq[ǰ�nt)�諴�����;UJY 6�R�F�D�|����{��/��<THA�"�������ҡNl��V&�ob��b"-S����񾕏��-=9�N'��|� �_�}?̲��v��d�`�I��K�GK�M���;T�C��OS��ʟ
͋��|r�&�6�/ݴFɇ�װ�jtj��-Q�mM��m~�J�a�����4�l^~�=�>R�����;��+KMC���!�Շ�vw���)�Z���)�xm^�M�~f�;yh��v���@5?�Y�����U:�uy��B��!&3m����l���U9�N�6�Ph�y��s:Ņ�x`�JhQ,I�Tx�`<��9�lB�&�Q%!3ݭ�V�:��
��`^�#%�����3Ȃ;?�׊�����$�b�h�m�bfc�:]5O*�(��L�X�NM�%�=�&GnI�����w������}�#��m��a�sbi�w�u�W��Z����j�{�������h����������Z�0�PH��hgz��������sW���� ���$�vE	�\��H�u��uʥ��N�d��3q�/Z6�.��z�3�+�k�qG��ȩ�){ �8���nJ�3E[��A���+L
���xM��;^虖С���i�h��О
���jL�������>W��x�ؕ��cS@��{Md�\h(-�ά�����e,t����7Z�������ݹ�/��h�?�ii�9]��J�M#��ePV��e������d�-X������A����&Si�M�΁h���'X���O�m��b����"��<����^���y{�y�il�H�_����SG&�Fj\P�B*�V���}�<���g��g��<n��Ƿ���2�-})�KG+F�;k��7��
�s�l?l��\	O�R�$V$�X������;:�l
YP8�fS�A])�i��T����,�����+#���lp`������$����鬦�]����l�z��g���ꪲ����
 o$o /2�y*7Y�x]D����|�(��-p.��X��#R�8�:�r��HUL~��%�(�UP�u"����ߕv���`�C�,�Q�`m	����ͅ^M�S<:n\~�w��z-@�}᫿m�i7���
}����!�]]��f��Д,��E�m}O�^��GX٦����;�A3T�ĄYQ�K6J�J|��I1z0߁H�:n���y�ek��b��b�b�����Mq�����&��W$�����1�����/��)`�fߓb�ͣ��Pv�!<�>�����Ċ᷸N���[�b��D*y����n��BF7�"OZ5 b� &;�ē*����GǬ���(H0��#�"��ں��Y�_��֏�B��+��|#�B�R~U���cU��R2iT��Y5*Y0*�1*�1*�k�o��Z�Yĭ��
Y~�>ia�!�׌Q��V���[�[�5XG��#<%�ͤ�;eX�����ݺ�7:��uU��p�p�°��z�~���d������͑��m��{r{EE�ͿA���q�&p��)Q�0?\��~����P~�|u)�ٕ�5.��B���XKb�4$u��'�j�ec�K�V]O�{��Ejܨ�2���j`~���j��E�d 2SZfbp�n��F73j)�O��{�.�%7q���I�@�أ��������]bKè:jh/����z��)�Tm���6��gZy�W�-���>|+�^S�C�"���娄3�V����}0����n�g��a5�� �K�K=XJ���#�)o"R�����W�?�ȝ	�$z��6Y����tzQ���/U��K\�h�7w��'��K�DlFu:�s��8����
��?NS!����z��~�6�M4yX��:��3�YfZ$���/�y�E��J�Э�%0^���jdnX�VY{���rO��O`�{֕U�qq����&����ڢ��OSL�=���1�}�������As�E7i�1�W&=Y]��XB3�*b
Ҍ*f��D������^p�.��n�c�*��>I��y��y��*�T
�U/��(�mCEC�l��F7m������:]v0Y���G�Q<}�R/�d}�:w�������f�,]e�Ft��j7���������)�(|�7vJ�������j3����M�M��7˞�������d�r���{m<�W����<�LɅRq��`�k�S�N�@�W��=N�����t��~\É�68z���#5~�lm�w���CL�8������D�Tڜi�~�"�#�,��IV4�`E}��U���a]=�L�Z����Z��)��Y,���һ�#XJzG�=RK�)�����2�i:e�v��E�H�W���7yc�Y���^S��"iYE���m�R�۩5~=\q�1�!�ưT����;=��swr��Zb�OF���%���4 �Ҿ|�)���4N+��G�'ણ���E���ƛo���v��vlX�:��4��B+�,Y;���Ϝ�HT[�����"�ؚ����1
�X�D%\�������f��y>eE�U��[p��Yzx\�k뷕J�2��5�Y�.�h�I%(��R��6<�,�luuu������ޏ�e{$�r�����-+Q��������s~|���(Ξ�����nf�a�/&��BZ�H	،�Ry���d�x�%��fU,���m�:b?��z*���"�+�p`�
��9�>��"��օ��� ��^���T�J�f�h��);l�������8���Y�X��׊	����C˹��&�����nE
���cZ.�S�	xS���N	%�H���L�Y�m�X����7����
��j����M�o�ڙ`�gh��H��{��P���ao��d�R8ϡ�s�	�ۅ�5k{�����|�1����Iӿ�<��W��3��Ο3O|�&4�#4/�;|�S9G�1Hx07�q��5¸od^���θ?������f����R'&�b饒%Õ55}�?'.�>��L�cH\��
#��gDd����?Mm������X��#���L��]��myJvF?�����s��	O-YH0�p��{��zY>?��	0�F�(���6�D�_�2���Pյ7����Q��/MM�b[k��۷�����Y�G�9ꠤ���*�0e PZ��!�6�P6g�-�}3�y+(�8>��wS�����Xcg��K�����qM}{��-z����)'q�� �q5�,���Q�20�taS�Î��H�-���R!� �Z���b���T3t�S/�)'3�d����F�vݟ��ޘ��E[6J�C�R�ceu�_��DL$�����.h��<��}�)%|�M��V�����.wI<:\"Ƣ��%��3��|\�X	j��W�ER3<��-�va7�w5�sb�y�֛�h��[Vɥ�z������L�f��3��mkiZ����&#D�x6����J��/�a`!��ª��_N�Q!nS�ouGǺ����>�,�J0���?���Q|���ױ
��D��$��t�|��5F��A���ǿcxqOBr��ͩ��u�v��KV���c]{�V�����h��(Ş��:���T��
��%r��d�U �����Ps�6����ԃs%]�"�Y|��%��2���[Հ��<J(=.9��]���Ip����!��Z�.�	Q	�h~T�ZO���MZf�G����Kň���ǟ�|�TL� MPofn���h�q��͵񯌓��:�ｽ �٠�D�����������O��ƃ~���F)ǿ�� }���w�{���T$����n��Zv�΃�:�WWE[�Z�O�k�Z{N�ȑ}�����!�����Q�&m����j:U8L����
��뛚��Lр�p2��]os�(���}||���k:j�n3\�Xq��ǠNU� ��yd�L}|��Wa:ܧ����0��'��$`Y�ϵ��}���-�zbZ����W�z�ѵ���?��g;�ώS�H�}Q�u�s����# fUT(�L)�NX�$���Rg���{2[
Iijk�݇�`�h��O�	~�=Տ]�ܵ�k�e�ݕޗ�P)i7�^���(�,�e�Ǧ&+Z�s�c��q��8	��B��%�4���14�t+B6�j�&l�C�è�!2*��:̩��d9���%k{���#����ä�1�X>��˾gt����}��s	b�GV��Q���9��9vmnz, `¬���՟z`�G��¢��:����]��wv�����'�"���(�p��m`�W}��Џ{��o��R���	�;�)�U~�{ �@�}��ω�M�$E[�o^i��Oh�F�S����������%ֹor�Mx_�g.ï>��ȯnn����>M�w�.0�� �%�/mWcѽ�������� j���Y2�yf�K��h#9|�j�G��G����U*����.~9���0�X��D!�%������=tiZ��~�-}rpׯd����C�}�(Z���C���;f�E_@%r��r.1������*�$�����*~���}���fo�3 ��Vo�49�/ڃ]o�]��+�H�<���+TJ
���.�/8N�5��6h8�6%�P?IYaYdg��oU>g��E?ks��F�� ���3�;��8`�#?���g�H���{�c�?AqG��(���	r�P���ĐD�H�Z�!½�7��)]���վ���G%�����J0`P���ʱ�)��)}P���^I2ڸe��\���t���:=�!7��Ę\Լ �(���c?�>�'��l���/ �/�/tY���0���gV\�ϐH�r��)m<�/X}P�E���>ێ6�5�ɒ�E9��-�t� O�J��ť $Y̧z!��Nu߫�S�rz�ͨZ��]^�V<��_��k�=1dd���KK�E��d+M��M�Qf��M�H��])�䫪�C����@T�zɩ�g��(�2� ����������T��[��Bi��2�ͽՈ�n��B�M���K[$�t��؎1%����k^�K�s������%3��~�؜�t������cYm�2D�y�^?���+�
 ��A㞠󡾔���b��9&��{!-	�������n����U�k���-�[��� �M�@b�*7�����;;��<���+��R*U:]�j	$"ݛ쇪i��"l��t��8����M9�t���M��2 }*�rCbV�w�]�_^D��[��8g��|0Z�⻑́(��MaA���6�����!n]D�(��}�h��R�pJ��"eȕsww'8���Z?iQ-ܿ����19�����Ua�0�?��{@�x���W����2S<�Ú�=�NN��
�3�KX`#�.hv��Yy�T�%r�8 �w10ڻV-8�44@��E�5�da����=o���_5��G9TF
g�V��9�U߫������mz1+k���@ ����7>>t����^r(y@�/6��ʇ��_�~t�O�6�g�g�kr\���{�b�sg@O5��ƹ7�|P���ˣ��)����h�������[^·���;��c�{<=U5ͯ����2�1T�t��=�9շ�)��[�0����z��6���#�Eڂ���a`!���y���y��dp&!��0��!����@4�:��!�B�����c\ʎ��#t�:E��O�+�ECC��4��� ����0�[������ͭ����J?taܿ/����I`�C'N�<�l�hd�{������Ԁ�"�D�p�Kȍ�5����S�k�~Ԅ��~U޻]赔q��wǵ��ج�������,ll�U1k������4
7��(^6(�����NH��֗[x��s�3�P�:��^쯯�5��V﮴����9u@���=�F����@�K�z�:�hc ǳ�DM�<t~}���toZ����x྽�����ݝ6����i�μ���Df�����ݮ�����R�n�ոx$�F���x�W*�"�r�̈��m������������淅X͠/�������am�d��[�݊�E"��?v89��`w�:!Ynq��I����������Z�%�Z�^�J���/��7��ur����`8'�>����?(�IE�2��"T(��4�7Z�ˍ����ʎSC�*��.h��a^M��t�Nn��ǉ�0D���۾�7�������jd���ٳz���M��;�����N�\�{@70�����Lt����b̦q,2Lí����A��X&�
�J��ij��v�j1��2��w���@��n	�`�h���{ecY��6nΆ'��*��`n���:�d>�/��.���"�PmW�����ؖ'�a�[*~����۹ƞ�w-{Ч=1��I�^��²�6�:%��S���}��+��?�R�96���vO���f��,�-�+1�!t{�D3���z�w� M{�1y��>�'��￣���4����.*�M�ˇo���32Y[��5�`�19ߢx�XkLN��m��}}�{��Y���y��ݯ��d"�Eؽ�n��b�0�֯��M�6|�� �r���:�+[!�ЫrƱW����=>>9�y='{9�y�u��,�a츩z���6;��Q��
Go8ܽ���Wt>(��:uȩ��>����v�0?�9��]���W�(r���6EZ���8��/\|�x}>��;�Y��y��������)�`YPWl����ڣ��:�K�ݪO�ov� �� ��^jAP��l]"���\v�\�Ƹ�����K�g_iFO������`��k����y���.�G���$�W�� ltt�f�jeoK4 H����%�5��
�ܕ\V���j�P�k�|Sx0<ɤ`�3���[�ǪW�����ui��s��{�����k{��Lʃ��l��u�wv3��F��{��H�S�`�����H�xݏh˗������E�����5����x�;��=�k���k���-�n�|���&ƻ]�~�-�L:�ϑt�
�z��
�����,	����T���g�w�0�x��Un-�ؿ'���/���njεxC����XX(�C�V�檍�+�}S��ߗ����g*t[\wP��Lv�R�߀+�mol���vW�Wɦ���f��x�΀�E�j���R�����u�xfD���z�����1к�W�]�x�6CK��n����!�ú���i�&���D���-��Oi�FV^������<�FF;�;o?�+ȇ*6��Vv�R��|����-\r�+r��5��aJ����< 6���6�f\����CV�eZ����/j�mZ[��n��U�?46�?��P��"��U�/���Q��&'��N��o¶�9aL[��z�y<��}�^j�P�	zU�����Z���]��~�g�nW��V[.�޸q�����
��КS�pl���		��[�Y��#sl�����j{�Y6Z˟;*���|�~>��	��W���f	ǌ~~whs����o�/�_��PU�o�@�SMdo��h�WX�����L�_��>���֑�{�?Z�=;��]:u�d�ȷ~��-�y�gR��[WJV��l���@E+�jN|o��&2VX_B^��$ȸt�q�q�N8�/�E���џ�+��?��o���Mf�F��g���^1������n���2�k�U�|�#�i2����6h�������=lȌ���4-���������r$�Z�K�O�OG�q�̬U��z��4.�����k$�҉V��vsq'�^v���}1B��J�������\%���|�5���ڿ��Bt�4��Y޳�^y�B��CKp�+tP����s_�]��5BZ8$r�	�a؏@P���F���IlNmLeQ����D(΍�(���Ҕ'��
�QhD+�) Min�vT���F����X��r��_������ %��dT�|ԡ:������9Z04"l����Q�>��5�)w���$"UAF=a�|���"�����6��;�)��a�? G�&dr�����q˰K1�����^���M�d";P-�?�J�z\ж���oA�=ӈ] I�n	d�p�������5;�x�Ә�TMue�Yr3�U��������~�|o �)�Q�ׅuㅎd���zΊ��ˡ�dTŉ�'�_�)�Nc���n1�����mr�ޫ���^DT�ssۛ���� �?�`�4jL�nI��+o�����*5�V*['�<�q�Q,ka1�����A֪8�_ @n�p�Y�XU�eM�QT��9)ݙґ�����6�@�m�{�+B��jm*4��L��6��Z5�!�d9�}��I�'Փ�1WZ[4�	
T	YGY��%Y�zd��d�ER�Q�eJ_��ô�Sk�����?������6U�h������S�kP/>�a�� �3A�R�`���AX��8��=�XD��#V��c��~:���d̩&�2���;���r	_xcd*��$�#~C��϶gܝg�+�(��}2�EF��$��!��7}����Y��_n�n�hE��u��撯f�]�rV�������Z%pQa�h����)�>6z��F.k��b���:�~b����{l���<W�jv�o���*ɪP1M7|Hc�1�L����i��$����ص�i��Ƨ]�]�<g�t��=W���M�sG��;��������UQc�S��Y�ֆ,V!7��>��DZ�/K�HR�[��%b�\���}����k�r��0H�X���H~����o��,�I�[�G�wߵ�%v�ݵ�n`���Y�~�����X���;[��rv|\S�Կz�֊wvV/6���rx�}��}��Dz�x����C�ܕ��<�ߩ
^+��� !�6��ݹf-B�;o�7Ս�E��~*��R܈������nau�R ����*X";�nTnjqJ�6��`�&�K��Wmc��� ���B��/�yI����, �9[�1`;T��w.P4�Ѹ��o-��Dp��)6�[���3��yX;��f���������b��o���WZ8m�J�#�P����6--�f?��=%�Gcܱ��`�LjW�����C,���u�
r�B���r�I�v��jy1�i�$"���2P���<~�e��U��m��a-�>�j|��6ͤ�q
*�z�b�6�Lc�K��0���
e�*���~)H��{{�K�H�I���s�/mԄ�L��Ӌ��y��΃�����}Oh�c/#+�ܱ�z#�@����cp����T����ׇ�%�t����ɩ��}xwl����ex�7�b���OxΉ���|�	n��}Fv��ߤ���FE3�I{���:��u�;u�w9Ʒ���[H-D�ݝ�55����<�k�D����xA{���Ϸ�wD���zl39&	.ll5�5�+�������[{�����Z��H�|q��P��Nv��4/������������o���O��Ħ���1t��㳷ײu�����·��Օ5�3P��j��7V2=���^��025�����������⢕�}xU����+(f�أ���֊��M���_c,m%�~�4@6�7C�����L�~��Ҫܞ��W�%'�k��o�j�́g��T�dr���q3n���z���)�p�*Iӥَ�IX�kIc	���:x������&zL�l~g��c�-!�����K�:9�\���@__���޴�����}�s�s����^�u^1ð�Pj	��I�(q�}p�3���*���⛒�����Q'��ח�{��Kd=s5-wpk]���h�����5W�	��tv��v��}y��'x�4��Ȓb�%ꖕ�a)f�8T�&��{�~�h]�0y]=s����O���z����$�����O3ُ�fS�qz��t��l��z��{��������7��4���wg���uN ������
נ��ӯ[��/�+b��д��5(�ˁ�s);���ُ-���������/N���cOb��b�Pz�S���;h���*sl�Z�^M�B���=�ṣ��e��海��#؍*�vxE���V�rv������a#��/��+T���+�o����HH�^H��͍���^��,��*�qG]t�,E��G�����H$D�]ǜ��k�-���.*�zUURxT%�;SCH{��K�08����ZnL���D��B�e4P�h?�+Yd���@X�^v�1.�)�F���J��9��vx�y�*����I c
sy��U���
ޢ{�h��,��i~�|==�I�.�!II���B	�/����1�5�Fð�ҏ9ɑ�B���'߻�cEمhS{�<cD�nQ�(���r,�[I��_��o�2>hY��M��M���v���g��':�jL�L�GX1BN�@%
Ƴ��%�x&�B��咽�C�Ћc��f�<���$1ő2��Y�tB����4Xr|ġ���?h� 1�l%ԢHg��Lt�'	���ٯ��lF۔�*T��0g��?�le��eh�?�QȚ��+�3�b~�'��y����R1��c����M�gۀW�7ės{��7j��,�91�����@���#����܄q��a���f"ٗ�f�������z��� !������z�
�֙�Y����\{0���o������a+�a�{{�y��/�fvʎǦi	H3��6V�MY��a�	��F#.��QA��\��A.o�x�=�>/���7��SHI�N'34iC�GO�B�k��1Kދ��vy���n^��ɴ��j�e3�o�6U�T6Cl�D�m�/�tq}-g�כ~�	�1s� ���	�ӧ�����831�;֠]�uݥ]d���'?��%x��AV��e�l��_�5�DJ�U,9V(������gT��yi�C��m2(Q�aH�O�M��~�Y|�J�����s�0�2�P�q�L��
ٌ��L�*e˘��b�#l�J+��)���u/\��S��KEB�!u	�{��Iص*/<Wj��᳀��e��Ǽ���_%sT��E�a��S?���>+�?q��;5)7�I@MӪ�Y5����Y	���gk� !��'�(��:p����K"� �2�p/��/}n_/�����6'�HZ!��s�0:��<(��H6���g2¥SL����f������`0:������O��q.&���EQ�C�Ɩ �D_�jĖn���������V���G�5�2���3qɀ�I!�@؟���[�2�L<�h�a��d�c7A5��#�<�g������,�E��h>��W]�It��X���D��z��?�v<�_��e���o�*׻]ec(��o_��و�҃�U=RGg��`_�S�V�$�����!$����Ii�?\>U�i�ur�
�7N�o$B{�v��0�2��~6hT�ޚ7�:b�B�?��TE�d��
�x6[�d+�2Ó+��̎!4�0�V���QiRk�����>�j+(>2i�j��#�~CF=#�ڀ`�l[�y�FQ~�Gq
Y��U**� ��4�(=)3%+@R@u�g���L��=NL-��,u�d�ךQ�jHK��#����<6��/b��n�Q�܄vu�2�9��ab}�l&��x?��'��O�}K�#��C�%RJ��v7n����%�Ӏx	?��c��0���֯3�S��
�9���_����	^皢��������Ț˂��]ƚI5/�qE���H���؂˚ݓ\r�:XvZ9�u�à�ϫ0��"�A�]���cX��6< �U�t>g.c�6<�/���7ܱN��k/'k�M�M��M�����r������qD_|k!���}����+�E���z��ҪX�~t��'8.`+�c�^ifQ[�jT!�E�Keժ�Yx�z%�4�����2a����Φ	*�5BH���zVgd�^���c����yaՇWX6q!��|����}�KC2e�.W�����:�@ak-�!5�3�N�7����*D+����g���e>�ߔ_�m48�mGI�jY���PLI�N��v9��#isN�P᳌� �"��C��P>�}�iPT�m�C
6OA>2ݭ��U�s�'�����<�fO��
���,1��f1?9���R5X��'��<)���3�Z&�<DFR���k?��,?E��ό�e�Qn�['�����:����N�WV��6c�F|�;�ؐ���`D->��C9�Ci�$���F���W���I2�4}{�l�j_K'ˬ��� *�8�3���Ư���a5d?�n���b-zE���p�����au�� ��L�����ރ&ePJ?���[Q�2�����޴lBF�]em�꒘p�H v�Lcj)R��V�ᢐ1rN��ܵ�6څ�Y�HU���G�����R�a,KN���j��޷����ٺ�!�J�w�0�&�$C6�3B騃wS�ת)�� +5_&L�ӡqy����.���y�Z�P,���sv@ٽc<Ma���������rJ��r���R�M��]E�W2v�2oS�|x?"��=�A�2��Kݐ�S=y�;����&)A/v6�E��rR<H2�\��k5��/C�$�?I�z����	iŔ���uz��#�M�A\|"cp���S����U���A�u3�f9�E���*��q�`�ͱm]qx� ���:�5�@});�)%�D^��\�`��$����%���FO&>���H�<�$��"#=
^����k��e�K���}��b*���qKZQʃe�<��
L`V�� [l�T�I�~���W�1�ʼPA�s�U]�	k�����?=.:��q����L`��3:�����6��T�� �?����d/������tٜ��y�}W�zG|.S�[������UM�x�gxdq�?4��[A�T0���r���#�QȲj�Xh�2 �������OX�a��{V������jc��?�% }UڔL���8�@���c��{�	�L}d��LD3)Gڢ��ɰ��_#SG��ri�Q��i���ӑ�ض>�������
Ĳ$5�k|�}�߿��� _Zj[i�:�f�rg��?�����6�W	?�=�<�wx>�I�.E�f���Q�N�U��;�צ��#�����]��9�������JM���9x�rcpR	�!g9Hۯ$W\�C�=sTh�ķd�rz����#�~��Ni�JK�ͬ}�~�?:>��"���3�u� �z��:�Q����"�
u{>���������n�oxbL�]���5Z^d����P�O�ZrЫZ����m�4�nߎ�U:��f�G�.~#�A�����e���&ٛ�sC�т�65�Oh �YT�8p3ИLs��x7x��j�V����IZL�ԡ�୉��E����9���t�(�A��V ���~��`��J`������mj�|�A�>!!��V_�f��P  W8�>A6�[��g�27�1�~���1^h��v�nz8 \��\�b�^	_�P�(��L�S㗷I\&����z8� "�i�
�[�w��%�+T%�4Sv��=��KuǄ�.a<q��Q�����We.u&OE���=���',�!��/,�(oc�)��nk� �=��(�o��U�n�P�*M�5���d�ks9`�Ltk��JK�ܱKT��S���cI�q��^��|�E�-���[��O�(U��N��1U��)�Y��z� ����\����ol?Q�;0��o���	摣<S�l�[����z���^)�Q�v�dȦ�ƌ:,*Tk ��U�6���_�B�F����j ;8X�i3A��'-˂&2G�wWl`�f��Pb�ۃ�<)�?#�wc��e�Ѷ��޽�4A���m$=��.���x���X+n΂��h̥	�ӎ�a�R�������v�����N�[E�b�v����ϓ���a�פ�>#3�}�l�#����9<dJc3*��K�A�/�.	+�a3n�,B���=H��S���$V�$�����jd�y,�i$dұ&��Z�Ց�4״.,ed�6)6	Ӌ�˕N��(��k48�(,��(xΦ)�jE@4��v|�<v���?=�����c��D�T @:ԍ��X��~�R��PE*2*rg� ��&T�5rb�lU�3��B�t;���	�At�s�t��)����~�Ә:ǣ�Q�F�W>E/���9L08�jÇ<_>�Қ o�}�s1̰��\��,$	�� \3�jX��K��,�&�S�R�yl�F���<3G��\k�qD&��l$�S�i�,c:+5 |!͊���������]��ԍ!A,A��u���M��6�ᐥ�l�-�K��ˎ��i��(�g�,g�!�g�˸�4�	�;����,��}�	1���H��v�iC��s��@�\��� _j�k��~iIkD�	��G"��4�w�ʗ��F]\�pVņf��?Dj3h��m!RW�.�~A�X+�FR�f��Y�Y��6���6��̰��cŏK'��}�3�N�˿*�(�֪���#�Vt�1�닷�X��$�������[Y~�I�֙����7�'��#�q�-��~9������y�Ӕ���W�����n��i��a���'?6��㕱����а�9��1w���o�����GU����;�f@���؏m;�3�ԟ�Z{��E���y���Uʖ-�s��waDi���$zFi#ڳ�����82�}`J��:���z�q�c��oG{b����ҕ�#A��?���,�,r,{a��x��E*�u�4ǧd���iD�&�[�o�I��~��K��t@��G�I6-c�ltq1�XU���eFo1m�'v6����SA�?���L]�ս������}P���o�We!��
1s��2Q��:S`BX���cT<�	�b9*-:�*OZ�N��ę����ɜ���ueD���q�θ�b9��32l$�����r�dEw*��F�ƭ
��1^bY
�Q�/��%�Nک��(�qcg�cx�n
Q��c���U��}��I4zŴ�j��$
g�O�V�F���@��D�m�p7�=��4��-T�?av�"���iB@��gP�Z����G��_����wU�5+���Fb�������T�c�LU�|��ߩ����v_,I��Y��1#��~��8�oܢР�Y�R�{fC��4�V���u�u�m0˨�=Qc�J�1ut'}�P�lN%x���������

�_�����/�fe�:$�5/�j7��.����&뀏R�)t�14U�V��t���T_��~�aǎa�L/���i�i��e�#�\��q�{�(�r]��Q�ų�f���R�?o�s`K�p���KI�e���f�Co�o��ܿoE�43�wM���l>L��D�,sKh�
�H�MK�0Z�M��N���3`�|,�ds�+>R ��ՍZ%��@T�.3������^��a?C�]y���؏j*��;�G�U��=�B�Rܡ�;��%A�{)n��Jq��Np�Ń{qw+�Px?�}�e2Of�ܻw�9wv�, ؙ��U��a������Go��=Ld����B-C3�O�R6�bƔ�3�L%5 �y�Ϲ�bm�����J��LIo��(雿Z�%X�kW���8����x:�f���}XAَ��JN�n�f�J�L#�qq�1�>G�_^u�.-�~G ��=��݀�J�%io{�x�rD]&kDv�l�Cӝ�qgi�� �{ʵ��s��}U��!)33?;:Ƅ�V6Jş�yB?��YPN(��f�L�,T��^v\7 ���K�dR�p<���-�5���DtvK�J@��Ҙ���hL�R�1��\y�$���-���q�*�(�
+���qP��%G|!�oK)p��=�B oM4�����S�Woa]|��3L��C�nͥL��BH	�>��(���X%%�&��;���q�������=�C�f�nS,�ѩ�����澑H
�)_C��i8�]��i���x�&ЙEKO&H��v�����m�F�{ܪ����}����2�O&��E\���?
v�}Kճ�[���3f��=����+�L�������3�_�p�uH��@�N��t D�JR:�tF$,���Ia�[||5p�H�ҥI�B;�,�Ro�?�O#��M^A)c�.��0Vކ�7�eK��>��+(�ԎˢW�4u�7�'^1j�u���<"�g2��R�>8�[���ك����MZt�	�BR��	)��B�%H��C9�į��oAf�������y����gW0RG��S��y�������[��O�oS	��|c���'�z C�h<F�+Q�!�l*������g
����Ld?�Z�3�x��/�3"�qv_drǙC����ܪ�f�Yz��ʹ��R�i&�wi=o\�FO(�Y���P��yiCd��>c V�B��d��2��K�@e��EZ"�S@˂>܀<��3�Wp�q����Ź> I!&�3wZ2;��Uc��د��]u���8T�$e����D�UW�M�4XkC,b���R2�_�I���\� K��[���;�O�uG�a$*e���O��{$��aBӭX)AT�j:f����{\�)��U������>��l�pO$9WyA_M�3�Iy�W�.��W΢4�/14�oi��[��!$>�������s�����~?��� �6�0��c�+Rq��`�z)%L/Q�P�'SdbqAw�{���/��/��{��/|�/�yo���(����1[���e�'тp��Q���b�ӡ�Ҽ� ��]��o�|Q��?)C2խWJ�"w�Ĕv��?�j0b����;
�C���yz���}�))t�ā`�! >&g�zI�%|x/���o���V9:aK��:�7�2��=�!��#��mS+@*f��%�ѻ4�(�\�r�1-��TN�3bL2fB]�SZ �����{o��v���#E���jZ� �0�E4%��5)���	���POI3�rN���qۈ���H�	R��ɀmO�@Y<?�䭨v���>��W�K��:�
�P�K���\��,��CE�B�oF���M����=�7���p��L^@�c\\ވ����<���,���r�����?���{�;���gtV�w��/)�(����7Ӵ�(�Lu��t�e�'Ř�(�5��Ԝ�S�Ŋ�"���1��e��L	'�]b�p\S*��aQ��T�A}0�A��ؚ���`d,Bu?��i�bӽ��@O���G�C]�u)a1>}��_�
P���{)v�ɺ,�I��dP�/�Q%��җ���]�ᇮT# C�w�/B b)�2~�Fb�cO���g�gTz?�.y����k��G}��#�?8Ҳ��������3|��r���8�FyksJSp��7�B�G"�[c�I�K�Ğ}�g�8ZŔ�+���E��A�y�����>�����w׶��,~���>��"6.<�{�Ӛ��+��Jg/D��`'p�e��B-	�B��36��du�ŧ���
+`�Q��ÿ���PmQ
��4�p�#�����]��5�#�+�S�8��Y�q�%,ФܰZ�e�_�c&���Nr9N�&�G���w�-�e3<f�`��k#�g&�Ǳ�B����ז���$)��)�в��E16�%�O�!27��D_�fM���bxj:�(Ruw8�=(g��UGoi+:�өJ;f��(i4�����9��J~j9�SO�K�X��j�ߵ�C0eRρ����10n�W��zK�`��ph4֪g<r(��� ��7�t�a�\:|c�o_]p���_���7�����B4�����Y�"K�Պ�� �;��E�R�^����@��eV�o���ʠ�h�h�`f��r0��_,S�!��[,Sȵ�V�	���iRb�P2�k}��wf��_��b�7�=�c8��[��w������Y� FY,��K)I����V�$��(��LY�5f㴖�����'��9�S'��r����R��3�ԝ�����F)
����_+׺�11�"Yw�!����Z�օ `��q/=� � ��XʴӚV�Wᰌ���t/E���{z�vIR��601M�7 �y���baa���5
u��oZ0\7�7K����ǿ�.n�I!�mJ7���������wm�#,��{}���5z��W��_�M�̂�clH��|��G�%9M|�OV��Ϳ=d���͍�+B뭯�?����
�0e�q�m���%w��>���W�Կ~ڻ���ʲ�6�0�Ϸ�bh�j��'+�}O?p������h�s��Ͽ+p�4��r{wK����",s���>i�k��y��p�������鰾y��V�n����m�b\����pT�� �ˤ���3�����Z*ן���a0��4����O�ķ�x�0������[>��*�A�]�����=zRO�������HBjؘŉh�u�x.�p�J�иJ���|�ˋX��F��fm3�C:��砣���/�B�Q�S���E���ъ�V��5�ʍք��`���"8����ή�mϺY��&��s���tHE��M
�Zjr����G�E}R����������28B2�Ӫ�+�����dz�U���b�_��c�~.Z��Hwb�C��?[[�n_����d*�	���#������-E��o��26̢�K{�ݶ�<!#�ls�\N�yW�VJ*�7#k �E�1���Cǔ׼��!�J4c-~��?DG�	���W��PU�g�T�����Ӽ�����(�A�CU��|j���o�;�٥�|>��[v�ӵ��&C�b�:���f7���Y"��4Bm�O����:V��v��O�w�D�a�ٍ~��u6̀�X��sF�9������:F����pJR-�ڥh�B.�4I5�ɼs]�����~+�q�<Ah�E�r�Vyީ�Gz�0����[R���O}��Fuxg�����pO�
ꮁ��jt��&P�GՉ�YW���*�=\iw����ƪ59t�H=�g)�<��$�E'�w�2>��k;�:��CHb�f�8��@.2�
{�(깔h���.��b�_���RKp�t��y0r[���u��1��~Tn{��` ��ԣ2;���[Z����}��MH�ܺ���H>��hw\���1�w��TƆY�Oͩ��(�rHXĘ�1/*�%bۯx���M�9[DBg�C�S���hI��AE��;�u�X���N
��`Y�A=�h�5��(�g��!�/��T/���8�G4fэЍOX#S1S4��$A�׈�QM'�It��.аі�n�ߋۯ7���"F��o���)�ezp�e�UM%�Pp��j�EK�%�v�����)oV�������NQ������QL�tx�ȼ���m�_��!���t�QH6|�F��R 
����Y��$C(>��7���v�HA���Ru�l��!�(�����>�}Y�6St��ٷ7���T���l"?/'F����=��ߴ~U�)}^gZ<*������b�a_�k��k?t�E�1$����(PT��1�Cb��3�0��?e��v�I,+F����w�1�)�{��C�mf�45��JY�1��X�F�21\D������Q���z:�|d#��
'���"Ō:J|M���������LR�ڋWs&׾�+����ﾭ�xfI��@E����*E�F� 陴�c�og�e��e�/[�s�v	��*��D�x�dy����*<�2����Bk��+�]K���Yl��$b^��r��K*E;6账}Y� �rEcW�C�FP�����H�tJ�ʐI�9;2�p��*�d����6C��,�ʃsR_�?�na��=�N�"=+\N�K,W$���¸�/��!�Y/i��MN�5h�g�G�I;I���`Ъ\:���f�5�4�k��՘�ig���5(�F]�'�Y�q�Al�A>�H-�yBS�P~2z�'��7�N�s`7eV�`�6T�����8��%,�^�lW5�ɥ7��� ����6.��Ya�<�x`.I Ր�6)�
93��#%�N).b5��5�:�/!�����:�EP)iI�}���i��Ӕ���;,~���8��)��:Ȫ@f3��1�V���$��&�1�	���/�Rr*UA4��[bk���r�����-���k��p���a���]��pa��T�?%����PU��ՀI�`�cZ
x��GI/H�䑠r
��u)��rM5�*&0?��М�,6EV���q�4��Mg ?ӷ���k���v�|���f���S:���d�����en)�F���3�D�f#E�#�=_Bi�t�(kN�I���fO_,2,�=cM1e�����ڐ��=3 �99!�7��TL�� ��3�s.��1�1 �Y ��Լ�G��r$Ê�᫢�����1����5��A�r�EbHp
��3�K0�q^�4o.jdd=�����*��,W�$��STC�������� mo;��p�T���Q�#�$E(4��4��QDlgP�S��g#+��W��P�f�JI$���M�B1�A�$v|�����?J9V����K����۵���_�_���z��Wg�
�;����;�K'�Ȭ�*�q�������F=s��nwRL%t�WY��VF9RZ ��pk��4��Zi�ʇ&5��	��]_g��.,EXlK'��O���^S7��kL4F��#���GO�, ���tC)*Oyɘ3U�F�2�G��´�(��$�v/\eF�5�����`F|��ʤi&�K��"ø��rô9Fx�SƠ�r�	�l��V)A�Ќ�\E����eҍ�d[���CE*vÍyRO'�on%���ؑϑBnXN$<�E����5�"��4�e�_�__l?�<�7-c$��Y�ِ�6�#H��K�ԍ��Mㅦ�ie�Ԛ��o��4��'q��/~qP���0�cv|��B���RH*�����̣��`ɜ�0�r��<�|�ʕK�����_��7�HD&�P?����fԲ��{}�@O��TM=h8y���cX������>H�L��J)���<݁�Q�x.b5LR?.]D���U����y2���~�\�/�����#>\d�3�ӄ�٦�g�������Vw����/<�<��L�I���e�W��/K���0�
��_Cm:�###��ֳ5I��E�;�Dn"����*z�a�JB}}���4���NݼU��֢}����$�4#�0��ɗ��L]?!�ݪ݁����P�|��#lx�g}lD=)t��4�C�5��9�i)�$F�i��B�j�MWY�w�����,s�{Jd��i���V{�D��iE�����I��٨�S���e������MMMD׏-ӊWڦI��Q�����whܴ�ܦ����k65(1Q3���_V���NQ[��;�E����HU!>~�]}�D�Yrw���������1�V
�+�W��(
wO�mR��yu��e3��r�c���E/���Q�����B3����GO���W!��v���4�<�g�@���;j��J��� �J�5H��i�E ��7��,	�K��hN!��Y&�?V��r�6!����)k�H�NV�zOT��*.�_��O��:}�$���&`hx۱���ͼ���7�6U�~,֏���S�]o q�n���U���k���v�Ҙ�^Ȑ���3Rm�lX0Q��Y���oS�.�J�u�cm��e���˗�^��-1��rv��2��,�,�mNq��٣.��_Qv�o7%�޽�2z�����y������	ڬ��&	e��.L�<�W����igR�/u5-B eZ��E�2���|؟p��Ad7]nZ����;n�f�۟%a*W������:�����o�?�jsx�&c*��rf���/���B�f�C�%F�,N2Ĭ;�Α����q�1��֌ꏟu��"��|�lXYݳgK u$̊�6CJ���!��@1�^�{cxM&��Om6u�[�t ��i�ZVT�g�b��Ѷ���*�!�/�}F�f�[\α�����-��FG�yG��Lx�@�n��[��x�Qc�៕�D��Rʹ=}�0VP��V�VQEݱ�-��
�{}��������\��w�}o��24V\è��J!
�V=�(q2t�#��KVm���`��v����;�c����bӆ�4����"�ʗ�G�+���J���/;3�Q�F����[����P���D���}UiB��4����������#�@}��!�� G>m�xqRe����<6<Y<Y��n�*��:�!ƕ�4_�7a��U���$q�zH��7�L �K�9+�i�[���#s=��_%�+�,]<�3�Hl\�d���5�=�
�2?�hd�dm��s|d����=#]�}�dżM��z� e����T�>�Ը����%��!�:Kp�:�jڧ���B��5	��������}�"QH
���e��̄���u�J�>�����>NuC����3X"Y�X�V6�ˑ߆�$f�쭑��jO����!�9��@�
Eݳ��E�Ø!`�'Q#o |BUi^�R�5c�}�g��_h��JlzG�z����(���Xr�=��W��5T�*;+��9>t��u�_�j.���_:��;��|~�
����0���9�d3�����D�XsMW��&��p(Jk����a�)�2>u�H�Aw�k[E̒x(��S�%:�+�F;�K�!$2���,4�|�����g�٘Z��'4��E}�$X�]�J�*���>m:JT.�k����+Jf�����#2D�tȕ�XX���������uH��(ԣ�`�a�V�@�Rh����_q���<*8���}Pg�eŭRV��z�Cs�@���˔>�q�	�Z���8d�>�EI Q�'�z`&Ku��ODEx���?R�~�N��O��}1��͑�뎾T~�}��\�b'�|=3:6�Ho���S[�j<Ԓ����;Q����4r��S�#ShR�.d�o��xت��V�8���<%ө1�8�z�]��n��[��+����u-�����gs�$J�AS�1�4 �" &\&��P���R�)�'���@x��#���c�MMo���{��{Ĺޏ6o�KK$���nH����\x
ŉ&���d�, �v�Uþ?PD�����	�ŕ�gr�'u��"~^K�vAI�U�8b��^��U[�<�G�pǕ}��Ž!�C�����mE���Ip,E�~�#i�/��3�����	LX�<��y��P�@�;��/�����q�h�(�	h������zz�GXF�ء��3 ���g?�F���Y�X�����n�D��iju�XuZ(>�"F�sR�'��h�����q���j��Sמ��M9�U[����laϸ�Y����i�x����Eh胷>��&-�R�KG���N?%y+1晆~#Nx�h(.Ҿ�֦��Уx�<L�OJb.��ud�v	j�Vwf����!�����:�vrh(�э�WQ��~9����+�k�ܑ�Cp����VR���j���)����x\�S|�'��#x+���V�Bw	ڢG�F���}:T<kG����'rJ�s Se��uEntޛ(?"���r���J�Q�����D�M
Lq&����X��]X1�E�^yB�Jx1�v��@��h�V��}C�o����-};�E�h���6��Z�@\�97��~ݔ-��q�Q��j孱��7�|#[�P���}m]R=@�7T��M�e�5>��c	�K�)����	�LVQ~����\��ק�L-�^Pl�V��pa����}���bg6�����{���~�V�^�w�T�R	���/Ag\��#�YY��\��_r,M H(�J���O<��C�~���Ϣ����ZR��| �,IV���Î���;sb�L)�
�ɴ
Tgii����U%�;e[���2򓽣���-[SS��O���$J�C��8��ǋH��NO自�꺟?%�V�G>�r׶��l�'�w��[-N`3L�����~M�U�qZ?�1h��u�m��]��)?�8���'�?=`_�-�)��ᏸ��~Ճ�B[����Q��m�G��/[k���v7!��]of�y�y����⁣���N�sB���+-��9�5k&�y�[�eU�?�û�Tug.ʠ��$j�$#��p�1�1�9p�*ぽ�tr�pO�c������%�g�m1\# �Z�lk6�>�^e⬭.��56��|1�4d5���K�Q��C�K.�޾Ziu5�p	���M�&d��Ɋ�Z��N�UM��M��c-�Z<l��h�j ��<���6���]�W��=���V�:<�-|�;:�;^ȃ��>�����`|���`���"����ۺ���<�W�.x��U�8	++�=\㺫g� om�/���ye�$��A&�b�w�=)��vt��QF(���В6Z��s��d��˿'��5A>�"Tq+ݐ�!��T�c���?rc�д�d��bZ\���_�o��
_c���m��XY��|��~Nq1g�OtNĆ�~��7�|��P�\��ˉJ_ej�,,Z��Ù�I;����k��x��L'�����ȋU�GR-	T�y@9p~�w���A%!�y���n�S$Zx-��9D��I�&����IT�}�Ε���]&}�"�K�W��GLbW���b=�D�$䈕*���b�ì��)�}9ð.�x�Qd�L��\�����|�=���̯N�������[�֦X3o&Bf��cǫ���꾯'�<�E�f
������W:e���-#bhfʱ �:��G�S/�[7%�i�pÙ��_y��h�ZY����ݟ�l��������	=\s�a�^j7�pLe���$�!�_����+�"�O�(����ۑwe%�s7��L=�7�����}��}c�?-��@ݮ/����h����WN�yպnY{[�W"O��~#_��[keuFU�]�@ZAt�`��k�9�s^�W�P�8����g�g��t�6e������C8P˫��w L.	�3O�7yƵ3rN]��="#_c``m�.>�ˇRB[L3�@QS�!����6ͯ�f��&r�0\�R:e�i�%�8�$R�Z�C��
c'�������l2��P��9�r����2�"k�>�R�N���&�yL8�^������	���ST�����=�ԛ	�A��|:�ݵ��7;��.�����ݖ���7�*�}भ����^e�(���m��F���X�G*�"SND��,��f�P�S�����zUa?�yz�������8����Ml��uxxpO`��R��<zKi��71�wh���t+�+R��Rms��Wq>���Y7s5{��+X��yrڗ�p�T����>�V�����Wz����2��<^��=]�(rW��E�N3�܌����1�!�L�A?�.��l&t[��p&���l^��Nw��o��22�=�m�o� G�c�
� ��L�O�6ң2 �~	�r�s�c,.�}u������FJz�V�g�A�&0�_b���+:k=���V��28�c�L8��4�"��[��uu4�l;m�lӨϣ϶'���B��mf���܄\/:TR-t���TcyB�#�x	,E�5�t��$��f�	-�"��?�`|�[5��@���hQ_C����K�Y��Ⱥ9U�d�oaEwoR�4g�]`���"= H���"~�}��O;;�)��)?�ٌ�tz\}=[0���ڝ�ݪ��k�K �C.��ʶ�­ �\���=�U,��Y�۷4��-�C��"+���_���]9�Ѩ{[�M�4>���겅 QrI��^��xR��^/�y�v����u�o
8��r��6JٽG�V%��&�P�b�$ĨvV����73_�N}�O(L���S�@z�e��K�|z��D�粎vL��wo��	3C�BFF^�훖�������<^����ؚ���,6Q<���o�[�UUU��M@n讅(a_0x3A��;t�IA����+�;@i�sXO�r�v\C�xՔ�Lh����ЊS�.S�i1�ugg�*�]�;�L��ٲ���o��c���r�)�{	�'��pi���WH_}�o�?	�q�|%�%�|���|�M�7�'�fa�J�Qnxf{>TE�׆�P���b=��}���^mX���ӥ�1�|�;5�)�yz��y���~@|�#�߂��|+������w�~{�/�n�:!%y��}�`�r2	��m"��\��.�P�81�Q&�nAh���hP��d"�W�쫀���=!JHhKه� @G��Dl�is�P��B��]=�n�_W�����:]����<i,���������ʕ'�mX=!�j�Z�	����՚/���z�,�>�|����^;t�	F��,v�꽗��k`�"4䐦]p��wr򍏟��TQ������|���ׯ?� ݧ�x���t��(2Ş1�f�V��
�fVE��� 973�GSҎl�5O�Fmmw#�[�F6$�v+:oӼ<ڨ�ZSe2����n����v����	�=�c��Zqg̗����CS�Tl��;�s#lc��xUza���z�[K���`o�&Z`�r��f�����L-ҹ�-�}�˧e�etyibe�_�\�b�Κ��Ǒ[�h'����T�7�
���q<�F-E풲�6�f�D�-|�f������8����"��lgd���@�A3�LP�F+�[�r��kIi+����:4+�A �0'�;��U(��3��Tz�`�?2x�V�vn�'O,����&�*���gc��1�h���l3+ϴ�1���V�'�F�����i�F��3ݖ�޹)	=���:�a�M���Q�0#�c<��"����5�E]�tr�M����2+���|�rS&��1�M{{
�0���������Ή�e�CL�L����Oy�����Lp]����˂�b�:����Ǽ��-������������SG��zQ�
X�XM]�4�mi�
��Y[�ܹq����gB���{̹�ΏD�*�Q�'�"��J��.Q�� �]&��n�i�"t�2�g}%�����J{`�i��ÆL0���u�;��r�T��!�4��Y�aW�<���-Syi��ê`�{;^> Ѿ٭����R�^)��f�¹�PCE�nM-*=@W_��U������� p����o��NO���a=�i�)��:�����R?�"�t���#i��L��L�o�;S��$�B�5S'�.'���۸`��ƫ<~e�*�#�["7a&��l�-&<$�mgu�Ckk� %r����>vM�#ƙ6�D[�5�9)k�$ZoOEt;�{c����{&bl�3���.A9d���4�5�D^�%R�+���w�O�i��<��ŧ�x;���f5G�B���Ǻ��T�%8�v\E��[1V���;�e����<�/�'X�r%e���-3�ަ�\�	�2�p)���>�;�\P$#��(w\&`�\�~_(A*�IKk�����3����*)6�#���Tʹ���X9�%��y�գ�5Ox��T�y��H��3�jt�~G�,����,�+�L�)�6iC#1�?&�.;��F�> IM�+�U"��	¢s�c3����wG�ƶ�=�4IqK/wO��%��/S��͟����)��I���ٱ�5g�`�mmn��ڸ"6�Nn{A�*P	ďr$�,�DP��ŉ���2�8g�e�R���?W�"$��#вb����~B�t_/B��K��Z�⣷��2�!O�gi�'Z"3��_�{>��7���a�p[5V��=|��?�i���PW�᝞P��ʞ�Umɀ��%�i�MG�YG
_3���W	����,A��E,��i�mܬ�,���+�ב%l��Ug����$1j��z�;����E��}���uM��)�7BM�ɣ�����⻏���UB9³F��[�#��݆��&�sښǦ��F����R�`ʁ�~�JO��{MA�n�kI�>A�F���{�#��*_��%G���[P�w
l�-�WO�YY�&���/E�^I�	��te�͏(���e�pN1�э�}�������l��m*ci;�DBnN��I�[M�\2�F�v��N��6���̂�����o���)KJZ��lao����鸠��'"o�)?�|���~�6��씖�ȪH�K�&`W�o��?�Χ�N�|ݸ���Q�K��)�!���l'u�E�	چ�,(����j������\���ƻ/����-�������hR��j��䶦a.eG�4湢��Fcf�u����yH�Xk�/��kR����7���;~�<���ص�|<�b*�3܉��6�tP�{����GM|1o������/�]Y�Q���*��%�&�.��L����t{{��������K����]g.B�I���6V���7=��aq��7�A�^��g�f��#�G$���-������f
M/1���8(�t�p�Ͽ���PB��������?�}���vс8�}��*S�v�4�zf���I�����v>��_�e9����U��=Ҳ����x����M��r�Ԩ�کn�#��D�F�uyXO�8w�H$�-GzD���Q/[���g�s�������F�#t��ֱG��8C=Ź��3@*�f�|�X�lauuJ��~���g1�TljE��b7*�J:E�4�����^1X'���K��a?e�_���cf~�V���PoBϽ.��'>�ť�W͝6�N�Pl#���P��V��G=��N?�U��ձ{付#��,�{=���G��d�@�){�HZRJ�i(��t��	[��Ҡ�`^<o���)�b	3�r�Y��a�7�Qc����H[ؕ����v/�I&$&���g���v��f"J �;��e�$Ҟ�:]l�V������ �	�O<�\�T�a��C��*>��z֬v��Y���ea�y�Gl����a1��i����s�?�k�E�;<��wC�L�3$'+;��܆ϱw���Bu�w��]c�P*�e�����ա���[�]
44����P��]�ľ�]h�i��ʂ��p�s���TG��@h���sZ
X�Z�ѢP"tL�f�܁]K�F7�f�Vս����	��=�W���
���sI%�9���+����XX6��
�țr��FC�@���R�7���hpJ�ۭ����|��^T�m�d�$�I�!xp���n�j���z��Fʿ��w��z$���.,"�(���?�Zy���_��r6P~n�'}���3y�����X�CS�L�;�������oGaB�����.l����Y M@���F��^)���1(��� /Z�X�Ѩ��N�����LuW�kr��
k`���?��f%�i��Q�V=U@��q3Q��D����0�r�s}}4�Mt+���(�V�'�x�t�J���Q�_,C�\'���e��k�5|<����O' ə��
I�-���q;V��G�8+����$U%�f�8P���mls"�� �yÅҮ�������
k A�NG�r����~Nܾ����]�E�-4�l8�����Y���������Q%:�
x��?J�X��m���n1r4>ȢM�m�ݾ��۫w.�slsgk��"����td3l��������kFQ�P6�YE���	�׾����C�,���̂�5P���~َ��G��m*LQGE����o���4�;mvK�}�a�A�~�hЃ���]cēD� ��B(c#�ę��+��嵽}��W*y�|c��E���>Hnw���g��MĐ���>C�����|� ts��F�~������{(�M=5���r&^��L��߻AtQozj���IM34��F�ˡR�4�۟�+5�<��S��5��2cU|���ŕ�ѧ��J���^@�ҋ�C�i�&��?jqk	������g�0:��S=�I�XE�nz�G�񤙨�J�g�mD�SgI�m�
��8��gaR��Im3��Y�jS%`�6dՆS�����(�e/k����m$��\j���ݿzzF���yS�RGǾJ�}��������w��n����w�lpj=�yH?N����I�t�6��� �?u��o�@�6��Vo,� ����A���y�!�HŜ��q�mE�~+��L�oƌ��>r��Y
m�^qQ�0 �R��=��~�83��G��B_#*%9�ΰ@#΍�+��R��A��:M֯�m���7>�m�i{�:Li���8�-�����M�I`�P�Z&����v���N`�t%���Z�c$�Qh���J�'�����u�d��?3�ߺ�9�<�L5�pi�PSh�3��:��=�X��npZ�NG:�>td�J�6�w#e %����e'F��&�vi�鸶35�?;�"�?_K�C]U	ot��56�t�
g��N�e�X{Ma�ˋ_��nb?��y|�.>p[�`���3DP�_>���h�P���9¦Ρ�
�7�
6�	�B�HYY�0bI��'ႏy�?�W�n?gۯʇ�OK��:���[5$�@ݸ��#G����4�@C��9VȝŬJ�|i-1�i*K�M�8�)�DW1Դ:�����e����p��Э���Å�cI�ay�w"[�,�0NP2�Ta��/O�x�E��+~h�˙r!y%k�O�Ã��O�'��㚉�����vS�rOD� `Z"6�t��O�v"l�qa?����F*�M(����P\�4�O��]�"��"F4�|R��7��Y�;��|����q�<��7+�����"44�P���9�U�޽���WW߬�����	�΋�ܝ-
�t�t�hS��W�OD�������O3r�#��d����-4s��G���Ӓ�v���تCՖ
S������8�k�lq,j#�p�d
�&J,Q�K�?��oq����҈\�H�����8�H��:^�n2���)�6Hҡ���NcM
aI�`�Me��D��S���= L=����鹏+��A��RfmڻYT�~�*Z7/�D̼*0��}�N�)�;���U��bg�@�RѼCx��& ���.u/��#����]�O�{�~��f!�4W�R�Ɇ�8�#�0|z�P�I���f�Zj��Gss���(����?B����cO{�	��t�UKg
��:U�o�I�x����y��7I<�.��O�C����>`������\Bؓ~�)�w�=$��(ff�����N��\'�ɯ?�\�W���@�t#���^��Yh饧x�ϑ����eQ*'��e�q�%%sX�*�"e�@�q�ʽ� ��#�i�e�fb��i�f/M��l��m͛4��O�aQ�>����	�kO�j��J������m�Gi�4�	����so7�q
�*b�����6���p��3�v��t^8)l~��8��,�Ե4^�P���TU����{���2����~h�8������XZZ�/�C���nh\�6��i@I���a�;D�w��x2�殑�Ie�:7������7�,�Y������1m=�ѕٓ$���I\~i�����6�7=D�8;Z�U�fe�΍�zӨdwǷe|[����� �`���������+���L"����k�5�����3N�3�&���3bJ��r����g���'ƭ3ÌA?�~���bge�aU#��p.�tĞo�s2�螫��F��Am}c���Y��ϓ��	$+A���Mvd��aup��i�[y��Ѓ�+ّ5�;�h�,&S4���/����Tv��%��e�<Q�\�'D	h(�#�n��t����u��F�.JeL���������`2+h��W�ʂm�/@�F�7��褒^��}z
�=����w\Cc_t��/]�U��O���	e�����)܌|C��?��2��f�~�@��ŭ�]����]J���������"�b�A+^�w�K�M������9sάL;�1n�JE�;j�@Mw��=�<��51%�"5%�����1�ܖ"�<�3�XJ�;x��9�y�/,��^���c 6��J��f!!/���f��ptP5-�w��-��do��C�s駵�o�,�T�N�ڨ@��O>��#��eEmu��a�-�������Mf�4��-E�g���6u��\�Q쮹�u��0���3K�b�C�;�y���.fvV��[s<��m2�f�o�����;�'�������-�"o��ee]�{���N*.���a�/�S�F�fi��\��7�,q�O����Mԃ�,<��|�����YL�� ܦ�ܯ��W)⣂ͅx]�ԡ�����_L�����2�&O?-wl���W�ˣ�f���=�<�-$�Gݦ�eא��z�a"5��\��ٿmj��`�	�i3?��'#�-"�B��]w&��y��ؿ7�r�W�
��5�۴�/,>�^�g$tڱf.)X���:���E;r���ױ�-��a�V�������#8vWW׿"���6�~�~m}7	v�A�|I-�/�%��9	6	�\m}��֕��Gڔ�ǆ����=X���4|w��,'y6$O�e�e������`��r�@��I�&�#����D��`eeՂ�s���//�˶TR�$��s�q�吲Ъ�j����WEW��U�K>�SJ�Y�tw�����q>��<��sU�XmY��o߂\�nh��]�:�n�DB�:�S����$Z�q_7a���`�H$r�:�i��r�Nc2oUj�8����	y�P>��N�A�40�,۾�"��H䧕�B�L�׋��J�8�Տ����s��OhJ�S�ݏ��<��W:����ir��ib��r;��z<��/&�p�	�|�v�����zXy�]+�U����?�c�������1�1�kO�i*���O���JL|S�Kl,A��x����>����[�].�8�s0��꒕�uĭ|j]�Jls}@��ɒ���O_ ؾ�g:�z��0L�A-�� ;j�%0_�攜�"�� $��Y����yY����X�Ay��.-_%-y�q3�SN���b�ÿ~���q�2{��+u�m^�z��x��';���|*w�w����~F�vy�&Ayi���b
�rr"��j���obr��^8Z����?û���d��u�7P���Ň dq͕����I%Y9��]�l+7��P�j7]򓝽oR�ğ9oڟ��Nv�#Lw�Q�X���X��1%y��aB�}K�T�����12J��#�(뤥ǒ;�#���vV���ia�(�Fj|*��dl�e�u~3�5���M�q���y��k-��L.�Ĭ\�[=�;�!�p�)���+�� g��(#'�fr �P��f8��#����|����U�Ǚg��'��YߣCLx��c�1��L!�)RI*�
<�(p��T4�'�XҜO��X5��Y����Y88���r��G9��W���^Jx�ߠ��nx��3�����߫4�e��x�zldD1��6yh?|"���Nd�6��ob�Ћ�liU f�,@~����%0oj��_���^je'�쁈q<*^�J���'�ǎ����U*��녕����D���MfEB����a�)�I�/��:����y]{*�g��������U�cQ�t�^��ߨ���8��9'z�3_��~[Yy}�����x|��-G[�h�-`%(�U!'3NF��K��|^�ZWW�a?���b��A<ok�V6:���̴t�@^6�PYQ��/,��ޡ燏�-V2i�PdC �[�Q^!�znk^|�B�~���eDTm��t�G�i�5�%%�6)���ТZ�*��Z���*��/�h�6�a-��}���w��pn�f�K����zn�����)"Qi���%��ⶸ1�vLϛ����@��[O�2N�r��C�0��i (��O�}�'�5߽�<�<�mت�=���U���Ū�����P?m���7B_�{auA' ��K��j@�:����q|�40����w����~�T��[�u,�,��ҵ�ϱo^?�(LW�o��2a�#S��ӧ�cf�[���u`]'�6�(r���֬-�����_���d �����.g	���BSRx�e��o������W�*������3D��_����'�F26��&�Uh�K�m3�=B,���i2���a�|����c�q$1��g���Ch�&�)���'���>�U?����|/"�HJ�_A��d*�g�d\��l��S��d��E��Ui�13	�rBK���Ik�Z�?����U�U��KHR*�JN�H���aFF)�����FY�q�OQQ��:���D�04�T4ԛ��s8w��4���CN�K���2\����%�r.I�zߦ���|�}��,�tc1)�؃�V��O�SS ��]b� mN�v@��f�6	�PbH1�9�mM���̥�b�%�'L�j1�X-]o�\�������5����]�������\��r�s�5��!ﯣ��ܤ���"�%�522q�� �L�l��T4[*�����<�Y���<{V}�B �,.ә�N	���� ����[�����6�I�2e��
�Eu�����\?��W�2Cd�B�JK%��@#��zb�5=�D�a��{*D�3��^.����>�	��F��{&�$����|P�R�ѱ�T�	�.�͜@T/��<�W�x�N�\����h*���:	m��'+���Q���:����eE�?k̿l�2L#�NX12��YHj<����Y\kg6���騙������;�WdQR/��yi����,�@F7��4o
��#��P�Fhi�26�7�?z�{���X�Mc�����mK)R��h��3�&]���$a�{��e�=EV��m�x��X8�5�ay[��c�3K� ��n�&D�h5����J��V�&��ֵ��ݚ;��T�Ŏ��� ��;�Q_
��.����-����kw��;f�0<���A�-[[W���3�K��>1qs2%xw�ժ��K[��`Z��M=75��̞z��ɰW.�&5��p��Δ��&�#��$��#���
Y��#<���>�ۺEQ�S��slI"�8��C�������|z��z�Z����^���'��L�OO֥�$�&���sxMQii�؞^��G��������NMW���D2&P�k�;Zcuv\�1J�J4~�v.m���֮���+���D��ߩSt�Y��
�#��y��߂&ǣ*��T� ��߿�/��ʉR���y��R)~��e�@C6�G���HL��$"kF���g�9����cf`�I���{3Xi��3�f�F2�{���D�ir��5�\G�wx�$�V!�?	"VI��5H��i/�%~��]�ҪR
r��?�[C��	NBF�I_�����)��%�(0Ѩ�h����`[7ɷ��xFU?�Gҵ�z"�S;q�)t,�Xƍ�ՠ%�-��o���$\Q$}��M��==�Ag ؟B�5�<��'���-�O����c�ty�����$�_�	|l����Jr[�lĄ���p擓L_��w$]��ȸaV����?z�Ɵ�@)�+��fIm
*��]U�s␹*ox�:su���E�1��$J1�}ʯ㨌ڣB�nYrkf{	u�{��&0�~̟�f[� ���1��<��9z�6T_�
$��3s2 ����?��^����+��l���b�D������)q�5�z��������^�P�9nNBp��!8z�o1@�5{��2ª�}і ����R�xǙ���䅓���{ aX7�\WP�e�e�K���Ђ�݂��S�<���\8�����B�gn_�Ma�8�ʉ�"�9n�x-�y�i��k&%%�Hj\ú�d�,4��ıDm!�f�`�?�u��R<[.o�"ۿ��j�2+�l�� �ɲ�w�B��E-"�����r�۬#�bM����t�Ă�Uҫ�]ERJ���-C$r���m���#ю��7������:�嗲kB(*զ�,�"֨�#��;�Gq�Y�!�|T9�Uc�t���x���4�$���CN�W�'^O� Im-k�:�B�gT�IR�{�T���0�%t��L`�Í����#��k�;������������������!�}C�����T�T�H���0�-1�D�/A��Y�-AV�aϏΆK��R��_�@�C���~bLTZ�����Ʀ�>�b]��#�x���7�/��W�]�KI�$�O�jPz%��'��,�J�c��>><�E��;�9A�H(8��I��(N���xs�z}�fmi)�~�7�����t϶햌f�X�%�ϔ����+��G��S�S��A	SZ�DV@�tpf$�o+�b�(�|2���6�J�o�CJP?N��k1�g��g�j��)�0�B�j�d.�Ud=!@s��$�Zf�PT�R�~�M��݄&��UA��X��[]�����ؖ&�|2��'I�*�����hG6I�-��C�Vq�M~�ڭ���dkR�
s��Z��j��'��
��W����UA�v!�ǁNuj���y_v�dS"�����;���/k�{�8�ަ��ŔFҩ���d��~�s0.J��O��݊�7E�^�?]�=-Q,��Rb_��^Z��rJX�?�X#@^����W��>����C��<�?ǟ9A�"I2SJh�c����>�OPz��{�--�./���#�飧�Ӱ�Se�����CyP���~�c+�UfGͦ�Pk��>�q���,h-J*�Q�:��>b����6�*`V�K�l���=�D�暴ݘM���h",R4-��� [te�0��H��_�5�r�w��J$&��r�}�*�ɵ��v����� T2��\9�Y��$ܩ;��9��N���<+]��vu��f/����8������������>~<"z�lU%V�q� J�@�)��m�z{'VW�,�ψמ���,�����w~����E��X�`�͚���Y��:��۞�̪|������$R�����NC���;��|TM�8�t�)c�~�p.Y?	���bGEP��ZG	]��!4G�%M��JA�~�=xKZ >\�%_���1�����������WJ�QW)7��Y ��J9��Q`�C�m�~I��"�@S"a&��J�:��<&���V�D�sؘ��m�׿d{�<h�=S˸�g.
n
L�����]B[���B&_Hr��f:�vY��\�}R�o���h+yA��ȣ�.v^trvﾅd��w��)�)���B ��Lx�/[��4��Bl�B����H��
�c��:xU0��.'�|"���Ԁ���E�>��5!�D=�wr{�|spt0I���P8����ܚt*=�@��f��cAP�1(h�\S�D��J`B�y��R��T������]�&0|����2�Ƨ�%k���V�Qeupuu��5ߴ��
���J��G7��=���G|�@-�v��!l"H�I�!X����N�!^�9S�Evyhh�#��D���M��˗]�I;�"��`�%��\�OH;ׅÒL�,� c8�+?����l;����|���w"���`��&Di �3��<���i9�aVH4w��������{(H�*�[�A�B�bn#b<G,�L}�"���X:-c�5�P0r6n8.�buwE�����_��/�Dx%Uڎ��E0k_g((��,,�ߌ��m�E�m�Fs>�fk�e�-�:��`0U��.�"z��o���)�p��]j���E���T���tۗFv�}
�:�a�����%�����������r�p�������65�0g����o��&V���5�2F�6�9�'������^s������9���H5��|B�7�:�ߔ/m����դ�]\g��-�~��0y8�y�w�bn)�0�1��x{���6W��s����(?����"m�-�M4/�G���R�ӧ^iX���ܬV�� ��N��N�R�� �E��>�3c����c��r����e�1��!b4�w^]�&�}~k��3M��e|s�#���n��^��#�<���u�eū�j���Y`fSBB���#�U)��b�A��:ɑ���4��!9r����_�0��zX�E���@9Ɦz:�%�G+��@���i�x�L0�A�_���Z�_�qm����t�<�b_]-��Y:9qj�;��t��{��5��z��0�P&��I����^�*Q�i���Z��X T1N).:Ȩu�ow��PT��)�x��뒠j	ƻ���bm��[{hm��R��=[*D�w�s-Y��K.h��;��Z3O��(�v1Ļ�a��3�\����(V(����� ����Mg��A�MT�Z������������f�zU�O%V𙲽�zKR
(kc-�������;_&�E0��8�Kz�[�'�ܖ�H�a~��ae��U�h=~���4Q�sv�ح����#�y�)�ߺ�@2:���zb����R�5U�(*ӓ�om��!TE��z6UKٝUU9Cod f�Y��319K�U��o�ۨ�C�Z��-�%n�����_W�?!�b�̊�'�]fwH��u�a�t�}�N���oioys���qM���������9��ߡ��a���i��5@����8�f^^�v�%x$��\(=�7�r���ꉥ��<W__��t�����ً�R��Z7���m5��\X}�8Á�Q�e�ڮ�T� 'CF��ovz�o��4oȟ��I�{��>�{6�f���f��3�q���[;�d"�XsK��y�
z=rNzhӞ12m��9�4��35�d�V�4y#�Jm �C�z%B櫚$(o�,��o0m�����g��~�<°��=N��?]P9o����Z�T���!h �?�����
�vN��w;d���4�{x�]�y̵���˭�p p~ay���Mi�&g�~l����;�7�4������Vs�s^�hjk��O�-Ra��I&��:���2xQ����b�I�����ǤZ�v%|�m^�v^����Q�똼�����>L��$�w����ݢп�[zV���%G��(;^z��-�n�j����Ab��{g�ߛ�ȍ��F���5M1��ёۀҖ��|n����ֶs��nL� ��n����*j���=�_������&Gֲ�}Ѱ��C/��@��sv�:e�e*S����k^�y�6�Jnd�} j*��̜c�,]�#Q3��3�tyWzr���A�l����8�U_��eXj�ذ�F:�����RLI�%�v�M�+B���櫈���,�Y�=�8���|Od�������<��HeHN�$�nJ�D��̋_�����I��	8�Ӯ���Y���>>�Zr:�뽲#�)���y�LZ]n+ "���)�d��(ŲAR�W��!q�"F��/&�Ԝ��I� YŘ��uq��_-�*񝖶$v~����%�'|]�`8���x�3���~�$yDS��ݣ���nk���4AQ4�$i�>����9�Y3�E[�OM�I��d^�q��@���+�ʊ��I�D�%g(�!��`�����s����3L��c�	��w�s�p��6s�*7/w�+�u�I�x[��h�d2>d���~	0	z�@y'D[Dx�?�@1o�����z��7M�F�`o���؅�κ����&�tc��d5|���/�����:
3���Qѣ�S��l�bT��'ڴ�����Q��Bp�4�Շ���]��v�-�G{px\/�U��'�D�|��<����߅��/�ѹ)�I<�u�/ �ޗ�z�Z����he�?����H��}��"ֈ�zo�� u�;���������	rK� >�9�ޑ��@����}���o�{��k=c��;�9%^��/X�/)�[����}�m���D�f.|#���X�i��SМ9A8iރ�m�69��)�_$�,x�k/�h}�u�X}#����s<�lj��$�"���e��^H�u���e�uh�2�Rl@*�J������u�/��N�f��to�T��N��6�P�ТP5��������_[=�޵2�LDs�g�;ip�h(�3Y��ݑi`:��Yr���r�+ڹ�A�;*F����7��$��$w�����V�X�}-��em�Ӱ��*���h�c]�9���G�kW�+���{�%�CB�`;&P=~z3P��o�M������q}$Spah�s�r�9���>����4r$X�$]�sƗ ����K�P��ܳ8x�I���i��X��ui3�S�F5�T �k^��R_[����dg�!�7w�=�%�޺�?���K�G�`�4=�>e/�oz5yQ{%�h,WO�d������@ #�o�4�I�����϶�~a����͛ �M��zOsz%���$!<��P6F���#l�ϯ�m� L�bOq����F�9~`@��\0위q�����o!��eoI�<�%� k��ãp��	�"�^�(VgN�a��8\@T��з�h�9'�w��y���1[#���ٶy�T?h���u�`�es����m�*�u��s���E�pz|5�'�׵!'<Q�}R��ț+�\�(���R���'��B�%|��Y>�dy�iz7�����Ą;O�}}�t]KLjX��$��敶9A�����3"^��3���:᱊ͼ��0�m���&Ï'o�3g\Õ�ok�>�"��8��n���{�	� ��[�$�v�|���ʯ�'��%���O����a�p�?d�@G=6A��Z�^F�e�n��6�"��n����8�U��sѩ wĩ�{�b-F�Ə��Щ�H~����U���榦�����#dv5����\$ػ�,�%ԏO�}�f\\���Ǆ~O;��Ǻ�wR�xS��`BNN���a��1�[�,��uj�z
NE��l����I���q�x{���7���)|j
Z �����Μ<�����n�:��0���t�:f!���	W����B�M��K8�3+LҔ�f�б��0�e~:Ք[��
�3��� ��	AQ�
�@��w����K��Q��7�Y��p��ĸ����V�;�&�k�Y�4Z�q�S�*;����_��#U[fW�1�p���7 ~�yE�L���� Ox��:�NKIl�r�����f�q���@J�H҂2WA��/d��'Eb�w�9�I���vW����5y<R���ߓ,����JE�` ��w
�e��F�w��hߦ�5�n�C��o������ �1�GK=�ö��rB�� � O�g�b��q7Q��j�}�a�17�q��2eQ~�c��x�~��N����Wӯ��#0[|)�I��ǃ��+z'.&fee���Hq���x7P������G�ں�'�:�8�)��4o)A���)d��˞��/�P�L�����#�*b�$fQ<��d����9�P^B�	�F;8�i5s����g�"�+ޕO3�/��ڏ����9�<�,�
eb7�i[�YǬqk�����Y�'�
kk^��� :��^����W��_�D�ڮV��XOG6W�
��BЧ��NY�Td�\�\7W�~�:�њQ��]���;Z �@��]ѱ)s�#[Y��,X'��Ӆ_@K��!#Uk|`ݕ]�x	��Tf��E�ԞbU��(x��>e.�B4'X�P\�_�y�6�]�%�s �3����G�%S��y�t��d0�R(��C��}0��CK�gRs������;�������J>��Ο
�+�ot&����55����߻�-\��aӌ��tq����e��UiC��Z��)+�@%O����̌�cg]�����eZ֝_���4ql\�ݹ����iy���88敔	�� tZ$h��5��M��Hj����uw��'
��k�E�?�
��<\��n�X{��m嵯���o{WG~�\�ۊ�ʧ�v֊M5������]���x~�;�<P���S�#�
�u�W����^�"/u��Ը $�8�.���jfc����e�V��G�NW��n��N����M����ʜ���_gJ��~�o���e#�ʓ�>�����%\9�諯g�9�(oϭ��q�z�S9 #sb�a�Ȋ@�Oؐl(�QlNR�ug�������Z��0��Ց���1�Ǿ~	��X�����\g_���B(]t�������S�ƾ���uĔ���a��O��\����Y�����Aּ�!+����a/Mf񤻃Wܹ�R��g|u����(IV_�.�.


6Z8\��]���xS՛	x��1V������oN�9�&&&���v�9�Ѩ7P��������"=	��h�Y�?p�K�M�)M���<�?H{��[�ķ���9�&�n����3�V��_��i�V�4�!��ɧ�?�Q����Mp�4�QV�ܕ�꒩D0�o���n������{Ye_Dx�%b|��,�0�JJ
�Y�ɬ��V����Y��,"�_4E���C��1�w�^e�ʷus���1:��]����I��Ajefl�7��Si�w�Y���[F��y��0cV�_e�������)))Oo`����9i32���2N�|կ���������4��-���@EE�`�1��u
�lv�׿5�N����)!M����D�?9Yi|9�ơ��
/T���T��*J��k=I6��eJ#[S���d���S#��`�`F�+��S�7�s\<|d������w�$��������N���12�ׯ� ���jͺ{��+Ea�����FT����~U1�+�a�DW U�t]]�����@_������S ��8g�/�?��Q�d� 
���j�6���`>�*?nB�O��:����̢���z\q���+r@�,���wvq�ݘ��ޢ0��
�	#.vr�SxT�\<]�[����ֹ��n���u�����M�<4���8�Q�׹l��޲��7aLB3}L����ؠ֠�~���4٦����V�4s���<���GZ?I�E����Qa�����1)�G�	�Q�=�`�[<G�\�G�m���o6L��D���Lك��HG�j����
��`/�)��K��ǖb�I*���c���|�/z����{h�Jц`��z[}���Qa�^�͑��7� f�Az�$�{�<�P��ad����9�#U�tsq�{i������02V|o���_�����7ruu����,0u������ĭ��0��]o�O碰��i�nn��QŨ�C�~���p�?~ͮ��3푍kb�%1���zk�~`=�����/��vj�J����E��]c3�����q�� |� &�Vw�c��뢠��^`��P˦Y�����R�����)#�Ne�^�����:�N�����bnm�������{,�c�舨��:����x'T��_[_���]̢Dh.[�u�����Sq�8n��G�y�#b��E��<��'SG�e������0���!N�J/��͇�r]�����WD,�&�d�4~�$Hin@I�9�[r_o�˫���0o%�ʩ��nq�Y1�_�
�|1��Z�?�C^��_'�V1[,򚚋7�}�W��n��àl�]�]���O�X5��Bl�(��B�bK5�,<C]��~"LT{K�;(u�n��N������vNG��xi�����2tu� �$ll���^>,-��A�}�9aa�G' 	f����7���������e�Ⲑ���(�o�^U��cmc���ł��߇� �a[����o^��?«w��q���J�I=]Ԡl���樳 ����-Z|���F(cv� ��M����ӂ���ڳXD�0A#(<ѽhaΠF����`B���)��-�}͗g�>�V���/�@wRv�l2 aҿ�K'ZѣSUU���\gqZ��j=�8EL[Ic�!���~�ݷw�N����Ş��
**�**�^S�T�>�.�b�Ȱ`L���A�M�d��JF"pJ>=��r��2���L��CT���[�}=����m֤Ǵ��P�i`�\M��{������xU�% �|\�L��L�{:5�M�Ͻ�����hצ~q�ǀ��é�k��ο�7/�/�t��c��34�F��
ŉ���$����������0/ƕ�I(O�36�t���tiiWM���C>퍒��5��f�eJj�2�c�Œ	�Y�<�����;p�U:��o��>��]7�Z�CO�Q�gA������zyVT�V��b�;�M�'��+!�p������b2�� u��б��3��{��ވ����:f�@�}8Og�"c�-5.V��]���ªxq�=O�N'9���j���Uђ�)���Z`&O��5�����-d���J��I\�f��~IeZ����{aa����a2K�>PB�}�yz���_#!%�G^c�~�/
k�Lx4)�UC��fR�*����s���KV��PbQ��c��C�N���]=��w��'�+�,D%B=�^���bp�=������މ�3|n����u��63'���ѫ�k�y�>APT�r��uv�{�ޢ(�㔊J���p�|E�ø��U���CX���@�,M��C�O�kӍ�����[gx�F���`h���CΕ�$�T�)X�X'���ҥ�(��3���Y����J"p���IyW�ye�~@>
~�D�p�`�v3I���-�=�(\_��h�wbn;�CZ������hԲ�şT�6>���+mn9�Å���!׫�Ue���ռ'����Al�O_Mo�L�q���6����퇉ɧ4 �����a���r
2}>Z���Ϛڎ���dS7������Z���&7����NFԪh�x���)��E0��9+a��D.Q��n%���1����Gd�cV����B.g=dYr��#&
_�+�k����ͅ�W.&`�<0�}\C��FT����a�ާ�S�S{�Hߚ�~��E��z��~��NY�����]3,�W:�	\{!tD1(E��Y
_����TG��l�ѿT$��<*2vu6���*��;%̛�9���^[��u���.kX^4i�䭔qyx��7�{��{�'�$�����0����S#�����g����ħ6YS�+��*�L����Q��9A�r�����e�{ߴ��%�U��x�gWCP�Ʀ���X���U2� �<ӭ�$���N>�{�-@�w���� ��d����}z�:^���/C�2���ݎ�^��4՜����u=~:����'|p|���>��/>><z	�Pg���2��k�J��ս�t��/"VB9��^��ܕ������b�^*��$j�4�9)���.,/���c����蠥�����$�d�d��x�S�̾��5ek���+6�7`��4:la��������C$�}_#�T��tv8��F�;/���E�����Lm�d��T�5�u�y	��x*���.�� of�������v����~/.ZY���QBt�������y:7��*��1���Jמ��)��qF�II�wΔ�G��W�>�_����>�fA�>�>�1XS��w��u�
�f.Uh�!� O(���a���-�#n�����u��+��y����m���k��K�i�<����Vݕ66���Ai?*jE_�v�W�xI�^��]���j�O
g��^on!3�{�����\�Ql�]Y�>W9��f����1VqSh$�ӿZ٫��v��u��r3����(z?m�2k��_������Y;��a��C�D�.oa��M2/2����sg_����G	�w	;�ݾ݁�CK�K7\������ǐ1���V>��r{q�����1������ yyU� b'�^{v�5�VF��HF�'2�G�%pJt�%�����B^��e_������f�3����2����d�<}!K�#��%I���h4Z�<6�`W�/އ�Q'��/KǞ�I��d��͖�ZB͖��_�1ӊ�2ݨǦ��h�^�É/!4\~����4�'m��w��1T*F�wㆸ�E�FJ�����6`v�,���)}l��-�6P�'O3��}���{}�}����q)�����78���9 �F]����������3�����14�H�@T��@E.��p�)I�o��/�$�#9��5Un�«w���d&*�-7y��x�#��`:��蒿��,�dZ;(�m���JiK�lr�HZ�d�0M_��3o9�>C��z  :'4��gՕƱ�g����O �꫘<7iī�zmN���72��d��9*�Dѐ3�5ƛ$h|
4O��"(Z�cL	2�����2�=2�t%z�wll/f�m�kM��;�Ŏ�t���;�:�'�*�7��h�������\��������<�Zm+���K�K��B���jׯ�k�W�O#���;m�������پ��m��Ê��F��M?k8���bՎ"8���9���)���ia�yY����YyVo�X\抰����g��V��9`|�+��"]	$�a�,������ēA��ދ�ݾ<^Ԑ�m�b��n~ۿ*�ÖE�/��3��P:�]�����y0���]!3���)�j �2pf�F�ܠyݰ_s���k�%�f�rť�Uc!X|�&,X�L��m>�{���_P�8C8�Y@TͮDH��.�pߞ*���G�t�?�:���E�Ԍ]5���ۭ��Er��=�珫><;tHCHj�5b�gj�o꺕�unZd�,��r�������#�5�y� �:��;�qU� ����,��<����|S.*��~7�e�+=;�E(D��{K�h�n���@���k�Ԭ�3���W!|w��a�of9����E�D�d�_����S����X�"�塟���������[<�u���p����z �������g�;P���QqH{�{h.8
O�}8��o����դ�Q#G:�Ά��0����a�2�nc���\�H��ki�,�ĒC��
'pڪ"��D*5�$��&��sz��$#Ń�"
���}��SmX:l��W�8��^�@����,�
֭����ME�y���\B���O�ax������
�%��������bu�C맻=���*2���"%0el�C_�C�.)���H�:��>��}����Z�#{��hoQ8�k1�E�n��Q�J?n3�:��;�=J �mX���ֿ=j�3/�F�8���U�'�5�ɦU%x�,��f����G�� ��Y�D��A�s#v�� �x�-��!<$j^=]�B�"����>dKr=�\?vH�+2�0������r쳳���R�T4�\�
����;RB�c�Ua�u.�Fd|�4���xF{tJ?AO�J��ځ�H���u^'����i�$������Yn����	`�>Y���~jg��:���^��o����vO�|����L�5�r�i���I�J��T���>��A<��[�`v�s��<�傿�i��3p�� �&�02:�����V3B�@c�w�u������
5��JEW���˘��_�ߛrh��=�xn��+5ɑ2����.�Gk��jp[M��5��eb��u�{a���ku��f6���`�=\�wr���d���!j��ζ3��J��k�o���U+Ơ<{2JͲ�g?Q_�0Ts��$�djY�ɟ8���v�E���V��i��T�b�[2��v��e֙��v8�&y�4�#25�
�q��'��\&	RqzLH��#�%�rP���{�lK���WY��%$`Y^�G���>3����zf{���K�;�����T�on��y-z�l%J��u9�=�Kٗ��1M]]IE��#H��+dٽ��y%�+�U�=܉��
�:��e�J�Lְ��S���������%�`�X��C-\�DP����g�Z������$<��p�%�`�����}�g�i�9�"#f�td�
���u/�	-gKt�SW���W��?�҇T��`�K�|�	*\�'�>�dbQ�L�-�+b��~,�?�k�Z��D�D���b4�D��ܫ��mCEbW��yr��D�Pf������>$�/_��a���T�ãU��� �8�wc��GٰͧIΰ�vo��T_&�����~���2�+M��Ӹ�Q�5���Ȑ+E �3U�'��^�0�P�Ќ�zۍ��8z��0�^�WaT�O�=�4Ѕ<����ӌu�{�������]�["l�ej9�[bK6h�u5%���?J$��"�q|�!�2��ف.���s_0BIl�%�����w���ރUD�h�ʝ$�)����� :;�)��D<�;3���儁k�mffd���ؓR[�w��b��d�cȉ��O�����<�w��z���^9F��y�%��j�M*�,:�Ш�g3�N��A5�3�Xz��"�c�S���3�����a�9:J�:���*�o(Y�{����.�ب:���e]�����Wf!�6�cm��`)�?��2(�f�~I�ww�,����%@����;,�[da��8A��#�j��LM���+�L_����)A�����9�@�z�D�o���L1�����tX�be��|��y�S����][qn����9+�/����tIf���5-��;�]�\�צ~O�!��Y�zOҺ'c��Ԍ4�v��ԕ�!����q�w���V2t����,0�?"mί��`��H|�����|b��އ
��t�-mXXk�u��Q��>|��Pį�薛&�~����Q��[~D5V��Vz5�5�bB���ws�ʞ�[5�"�(�J�rk.OG�����w>��Q����YzA�����k�j_&%R�ꃄ�IB.������,���|7��R�������
�`nts��~�A�Q���W�m�HL�p"v5�4g�K/]g���0���kC�$/�Wm
�.���*�`������d�e}�$*Y�S/k�P#�ܳ��g����w�`
܎� �鬧MƧ0�M�/9�/�<��r�@��M nN9��?�$�a����P��h}t��5���ċP��E�<3ǋ�����]r���o��u�$G2�n�Q������i���s�_��2W�s�����3��ο��G�]t��CHː��sUl�Ѭ�n��X���a�S�W�I���	���6W|E3ϟ=��'Nv�c
(��mP��w|��ɏ�L�Y�.�h9��̎_�M�JZ6���ZM���fA��G��qq�����$�'�Պg��^��;�j����x�n��2��E9���[������pK�A#�V�ܿ��04"?�|���rw���G���@��LDĳ����y�5�4v�]�˶.%�y����5Os�>�g�/D!�'\^��gla��_
�$K��;+3N z�Y��`e����/�˷�e	Ѹ�4b�N�R�K��S|��[����f?Fnjt29O�bǉ��n e2�e���>��7"�2�$����x�CP���b�pWYv\It;��4���/��I�]�m+[�]SV�o�"��.���k#�'�k��>{18��b�U��4E�{)Q1�^�v�V�iE%��:�vZ�|���3H� 8�MO]��{Zͻ���{��'+*F��E�UԐ�����4N��2������*�S�؊���.� I��N�A�i$1�;(���n�b��(?\�'%�$�/��-OAպ��Ј0_꧆
;���Uy��>�O��㊷�1/��dwfK�����=һ�x��^z��cͺ�9([��������U_��t�3[o�hE$*��Bӥ�����*[��Ҷ��K�F~u����N�j��ͥ�-z�2Nv\��s͑�q�N������TP��a�X�!��tBD:��
�m!&T%>���k����� ���k��g\>��AL�*�2�'ǩE'!4��;�XcmU�P��`b��@��u��Ѡ=v|�1�u��|�c������ ���O?*�L��N��Fx7�\~[:8�5`(�W����2n����n�=�e+ʄ��A0E�J��T���]v8?7H�W�l;EP5ݽ��^){��4x��;_X����I�IY*r:h�K++�Aa[���8��/5��:S�-�����\�ϸ�z����]&�i�j������VG����u�z�bъw8�U��U����g��V��A1c{8�>%<-�b�F&������������ FOOQ����+PۼGw ��Ntu��~M-�ڗY��T~��t��p	�kҴ�${<���b_Z�i��*7��d��}�'"�D������d�-qf��0������&Ժ@��P�+	��t42 �2w�ŌԩC|�b
�k���6���c>~U�4��.��8�D��%�Oɛж2Gy���Z{��l�hX���g�ҌJ��:��jš�a����ު��p�be��+�U�$.�zyI�<ϭ���8:8gAC�d�Sa�M]G�m���,?J}T-^���>���PY!D���dԠ��S ���xZ�x]aI��aQ� ���2��J#�ҲV	/#�/N].�MC�6^��X@b��u�����SѪ�ݦ����hI�G����y����px���q��DP �2*��4����������P���ѕqt���ޫ�G�U��+&���EԻ��6U��A�_M89;u�=3^�{tP*�,�"l9�
���a�A�^��ʙ<�gaS6�6Y=�m��6�^�;	wc��?�	�����^^���HTf]C�i��C��5pqK��=`�A0��p�|?0�a�#�<ca%W�N��:�e��΀��A{������!��������>������^I"����Yy9�ͺʩ�d��	��z�r�8#��n���{A�
�ܩS��f�r��h%J1�\�o��zY��4���113;�64�����n|YJ��^�`��
�+�e[�rl�C����O���h�5�P��ϩ[N��É� ���+OOYa��$A�Mz5`�u"�I/�-���a��%��h�2�=N�T�P2���v��^E�G7��H ʪ���!r/�XP2���Ǹ�.r^{�ǟ�M�����e~�������1��0�n�����PH������6/�3����А5�W������ZZ��j�	����]��Wך��1��Q��5q��4QLD{����k�_�:�%�OɫG/���h���d��c ���"j{Ab���&��ز'�^�E�\�+�i�'�}�����^�Cnn���c��D`������C�I9X�ŷ ��c9V�F�|_{��o0��d��0���p�F��]zu��n�I�C���k�������F�+��%�
�z}�n5&�C���@����I�ť��g��q�{�3F��\�J����Y���F����A"����&�]�?PF��N�{(�dJ�ر|�þ��p�m�D7{�J'��){wx/�.U��h�&8�10]��ׄ7��PP�?�$�����7�n��L�XêU������]}�/��u��Џ�撐���N���������ӘQn�}���b�Y��)䯙�$�A
���k_� ��$���B��P^���U�����?���+`0����)���'9�eH�����{>ҵ"��ZuPw���ڇ��8���ғ�V�7(7�-
�F6u�Y���<TUT�\^r^���5��`�q�X�o��d��%)�k٧��u?Z�6$�����P���Xi�3,��E�	���������=}�R$P�l���Y��s�p�V��;��.�9���9[��=��IU��"q�	�L]Aׂ3�EQ�"ɞ�B�1�8�\Wr���"\Zy���5^�!��̙3�Ɠ7`�[d��Y�@͑����-%؝��J�$�j9��cT��������_�vu1L��n��V~-b]��[m���\1�+��/�bE7�Z��E��"�u��!]=�[Y��S���`߸*�iA�����th��`�i �I�É��`��/}�xJ�F����v)�j�"���������_!�G�_?/P��L�y=̍ �Bg>��T_��?�CK󺏱-�.5ק�L�����.G}�(xb~�yx��x6�ܕ�d�v"VP�?b��S�j�Y_�n�%?����'�������#1q���/���7hb�4�-***X��剃�.�p4_�-��'�-��}P��\lk�j�m��133d���{M8�X��%�0>��}.�AR.�w��#�6Qn��*Tf}6	�i��3�5��9o��U��j�O(ں;�܁h�A�n��~}T�{�ss���*�||�k�9m��]𔹳����r����|N
��)�,����#�io_Z׳Ťʰ��%)p�q�0o�;`��
}��U����1�,�F���L�F�����Qjg���zu�h��,c���*Fj��3�?�"��(	��������Y���S��Fu�bԫ��}<u��gv����a�5���i��`po�,Pdl�4�G�I��%�+�w�s��	�v��K�ӟ��L�Q�ԩ^��R\	]�t�PNԋ|L+դ2��rJ�R���T�C��22�����d�b+R�Q�RG���R��A���}fY�\����ۤ�L�Y�*<V�M���W4 ���u7F>v�{�r'g��GMeu򘅸��������'D���!:����߇��Zz(U�Y?�0�fTD��CV�~��=��8�!F�	?lL����x����K�/�G�yx!�.Ol)��Ռ��8��3��;�u�8Ih���!� ���-���y%���	��/�p��k9�^�U_p_D�C.^����ę��4P�or���� �%>�l�VB��F
�k���9g� {�����G�@a��2����G�xx�:��6���U��?]s��2҆�f���!<����^����	o���c���\d�Lpb��z�����MUx�@u3�A��N�<� /
f>9aa΄;G�ǉ([�F�E�6�T���D!�J
��fN�?_�{^6߽Y^�SW���,�+)>���8���/�`.'��&sENh���A���c��,=I��w�d�Z��"�r�W��{�0+�Mf?�Q��H\��.;�>\2��k�e��Kf�l�p +�u�F;˕JP�֒��)���/�DR�l_g���Σ�$u���#ෆ�+EG�����r�h�b�8����j3��|k��=RK��y���2��~����T�� 3\I�D�?�e����>#8(:���-"�=+,�*) �p؉s���)���v���%�b�E���'�|<K���,:�0sH�\h���{�blӛ����)�����/|1i��Y��8��O*Pf`���R����1^XX����@X����	��2����΂��wyR��9::h�5N���C>�A<,��QG���� (�m�a�n�a�0����1=���K;���w�y���=p[xv,��d���H��eO��L*�[���cd]$�	�I�=nR��ץh���¡u���_�c�˱�p-�v�|%�izn8����ܤ�[��Q�si�@6y��I�U1���N�s6�j���=l���Js�h�KҤ���7�w8��cLKI���k�lrk�~n��U7�
G�d_���&�4[�N�9��#٪�a�=X�w�՗�j>�����F
���Z	�b1|��Q��\�]؊�:U���]^Z�/E=a*���ޒ�ɋ?�[��/$��s�J.��:����A���4�UW�t�㳼�V�x��G���P ����m���Z�`���	ŀ�|�0Cپ�#� Gz��i!�k�k���j�e[��pP�Sk�s1t�3�
w��R�_V0��1�,N�*�S a��߬��e�������5ϸ���p=l{/wRU����O�^9�]����e<fE�����x73�>���P��ۼT�T�J�;OX$�L+�laՆޱp�e�%��׬ulԼ}v'&PSR������]��3>��W�*Vl��?Y-%��bC|˹>��C&��]͂ A�
��*'��vOZLG�猱K�e��m�jh�~�1�B�	���=���a孶�!K�q���Gu��0�ڴC�8?�Յ��ařv��6��x��v�m��!W�ϏOq�/���>�)6"_�v����s3���4Ky;�A#�V��Cbͮ} �R��F�>~#�+G�O��lw����w�����/O��?Rc!kA�d���Fʧ����^��Hs�����J {?u�RĂ�O�Cz���������qs��]��ݻ�̖N�U��c��Ǌ�I{�F?c�H]���#��JDVj���F
ycF&F��U2�FH��8r��������k/�[��@�O�P(����ކ��g����q]|�����хa���Ps�����A�퉣��+��|ݚ��-8�W�;�>��Y̶�BCcG��8H�����R����{��T+r��ܼ�G��!�������,]�P�<LcG��J������777�<��x&at)c��8���]`
;7�\�uu��.z��r�Y�������@xL�Qt3��F��t�'�b�6e�8v`QC�%=&���[������,-�^��o��#�����Lw�S���T�M��3�"���h�����U���֫g���珟 ������6�EKv��)5�����zM��� L?�0�ԲAt}�6����!_���ǻ�j@+0�`/jÞB�j���A
s/��[U
c캩nm��C~���� �9���{#��w�U���E��n��:�D=�s�V\js�p�1L�Xy8.4�l]�j�����HM���,{<_
2���������_����/����k�2FJ��)E	oO��_ߐ0ɏ#��97���ߞ�~��~��&�o^Fq�OW�d�䯦���7�B�������$�]�~���*��fq{S뻺!{����/�Z5����Cqz�3�B��5�+��\+��E��n"���z$���QLMZ��aW<~�Ư�/O�4R�	�>��]��g��s:EZm�*'��]����,##C	�)A�:�1z��^�O��H�A�P�_�x��/a���l����-��Y�P��ڸ(g��9|�֯N]��WB���~HE'ݟ� �șj�n�dPP������λ��l�eP�����L������;xll3#��yXP�e�s��{\�W�3����n�xyyw{���r�q����B�ߞ��R���^�c*mc�S���lh�bk������R�z���h�p[��&�Xӿ�d1�d`���^3�x��jU�E񑿡�����9�8�	��-�y�o���?xFn�&��O4���z\W"144s�)�:��Y�=��r��F뼹�-���V8�U&�%_����,X���2������GR�#������vm������jQ��?�#H-���:;ɡ2���*��x�������ж���\�_S�����"'��3��0>�R�"c�8�m�ڨ���3ˮ0���9��$L�bB��ꎣ����Ğb(��bj���SM4�d��A�;pa�_�,<Cxy;BK�c!7�o"�%�X;B�J�Yq��`�%��g=�m�tV�a[�.c9H���g���= �9��w�������M��%dl0B�u���ݕR�_�Ȋ�K�_����Ð!�/� }R��12Ϧ���^s��b��>i�7��C��0l�u������U�i�_Pp�̵L��!�GĴ�&���I���]\��
׭�oh���< �����j��6�c(@x��5��3�F8�!�-���=�R���ʃ�y[ˠ�����O�u�&&���#cˌ)̉����TD�9�jb��'�NMi^�)H0[[22w߻��@�&и�Q�}�h�踆Yn?�h�_U�-�h�(6^��F��X2�Kt��>�-[�y��$�Y�Wo���u|+j��W]�97��;��D��3j�Q�Їb��ƌ�7�<���,�˖�SD�y@�dB���e��9�~]�/�7��w^���Wo�(�m��s�ф����%�g�g/��֊��:�i�=&p�R1v��C-�%�b����߇L&��oX��5����6x��`�Ѭ�"GK�.�*��H�t�.J��f#�ǐ�jv���WJ� ����\[.�k��,V�V�&g$��|�+��d�#����3����T�A?��П�����������B1pj:
%#A*�S���k��J�P3y����ka#��8s��V FN$���د��p�N]��ffIͩ��8u1���p<$z6��"�!W=��o_Cl�S�%�|��.��&�j%<&P�7�ws�^3YS��J���6�qN�Z�)���f^���7'�X[��7�2�L :$�#@E��a��,���A�.��K�����]tD�7n1Y|�`ۊ�R�ӏe����H#��Y�����w9��,e�܂f���B���o��ZF�M5�~���I�ֺ�;n�~�l���BW�}9�� ��:���cI4��~>��%�-�w5ڻf�R��Sq�C=ݿ���׌��"{''� �� ����5[����^ai��3G��
 K���o��.u��y亻qۈ�$c��:Pb��>pҽW!�wO�)ϭe�$��1�I�G�����ݽxJ<A���s��ވg��-����˷@.'������Ң��@��W�q����g_M�T���*5�����HSvC(�BJef��IBaE%�w�9-�a�X���T�4E���PNh��������8�Һ5�_˕31�U�{��pv9IVXp	���X��]Y�3V�c��t(��i��Jg�E��"���
݊;���������
�8��ş�_{T��;N��	R{�.�㮴�O'?g�`I��7���rq�*h4)Ѯ��������r7C���2c&r��_NN}����N�����r�DSlE!U9:���}&��-d�6_M�7w�j
(_Y	4�ŗLč��hN�8����*�g9��8R���{��g9�)��k��y,Jh���\ZӷQ�P'��uuuI��\0F������l_��%��
������7�L��u�v;�6���?�ɇ{�_@,��~nma��*] ��y� O���v�H�/�ylR o�!77���:�P��7�v�����s�����5��7D0Q��ٕ��<rq�,[Qad��9!F������x�M9��ς�IMf��
�C�l�I�y��A@&�4^�=�4�9k��G�L�\�G6��{
��;݊�W]���Y8A������#��>e߸dP%gD�3ᑣ5�s�v8)��Y�s��0�� *�q�>�D��I1�XPR	/e��?��E��s=�A�k/ʹ|d�&�4w��6+"u��y���h��_`��!T3��g�6���Bg[�~RY�_{v���i��}�0��OjA9�I��c���j�~q�3y�E!�m2�;@K=O�j�R"�Qׅ�d�$�P�Ok��vV# ��Q�>ϝn��-���?��	j����7^��%��_�r8�k�*{������%��f��g��/?�8�Y����P$+˅f�2H�	&4h	����e��پ��. bt4���sWnc�6�e�	�5��+��5��'�HX{6�..2Fk�n"�*`o|���n��e��R�m=��͑� �lb௖cM���to ��ހ�n�s8HơF빯����^$���{rv +����if����AZ"o�	���,4�O	g�;@���c6-v�lekia����ۛ�v���׸���?�lT����H
����JvЯ��e��,�QkU��3B���5Ⱦ�;�/�`7��NcU1��+B��[x��zX�q���V8PՎ�m�P^#U೹椊dW���<sL/���_�8ibl�5�����hW/������#\����o-D���$�ļ�Y��<p��������!�{@>LW�~�u�ʊ<#c��� 2]jX�=�@���8jb%j����������F���HV�K[���9�� �Ak�0S��ꒌ��v�OI�ZFG�m9�T�b��T��~'��N�"h�;�Od/�����۽6���V?-�nt��?���1�5DZ�{5�/Ʊ�W�l~#@u��\�7��	���?��&�_��I�J���0���k� �64x���kG��^\��CD'������J�~&�y��}��lk�qZ���γ����1s�������'��_E�����_D	iZ�;��H���n�,��-�3����ϟ�K��?�`��N��,����#�0<�u�
�S��Л�^�Q`�hR!zHƁ}�>F�m�lp��q�X�.�\�k��lW!E_��4�ǘ��c�����=O��(!��U�@�m��������|z%��<an��Â4v#R���'��{�َ�nei ��	���'�q�Vڵ������j+w��^arrM+��ogapO�/C�)����T��
.�2�Y�&�'@r��>��/��z�z(�����W����Y2xLD1F+�%��x��rV����ʜ�0]�{�K�Mj7���,��r�{��+)�T��IeI�r����:�%�[��,g���K;�F9��~��⟮����DVi7�הa0cp�p�6�����:�3�M�ӊ[;��?�,k3��-˙))�d��C)��|�Bۻ'�55��-���zԟ>���vܢ���t{���Dޞ���I��Κ;�v�_��ѱ��l���p��и��:}��>�xs�v�����٨i���y6m���R��\^�Q��0��j��}/
c�3�q�Z�(e�?�,ÜGh7�>��G����`�h��,�3��`�4^Μ�x-�
 ��c�^�g��=z���e�X���ƸC�����7?*�� t�øHt�M$��Α�,�0�����Cg� �R@�l.���Z{y��mŝ�%��,;[��Q<#Ek����"<иhW� ����)f�'�3�Q�G�u����!�tT�7��W�+hR���N�q�f+�^��u�ԥ��x����.�'x)@)�x[ �Y?�U�Cy\a�\R��8�oP�+��o���Ҝ�[�U�+���y���|t���K�^��|����T]`������(�ڤ���m#[F�zv���m9[�c�彇>��3�Q����G�c�)`"FA!*3���YVIn��IN`�w�;$�y�f�9.. -c��N�ʨ���f|F�>�Yag�A?��;}����<o�e2n�\o��hg�{g/"�>g��M��4�N�[��U�O�z J��6W�-"�7`�}��	d�V �y�Yk��wNirY��1�����Ϟm�q ��3�:^Mxak ��lr�ŝ��0�ї�j�����E=���_���kL��|G�� �6���DxŎL��ݤ���+�e"�
"+(ڠ"R[�+̲6�Ҁ�+��2�X�c�qJ��(EE���Ã\@آ!?y
�rGE�I�r�3�n<W��V�OJ*
6dA?��r�����u��Y|��'%~��`���,=����l���aLj�W%vwP�cE	Էg����}U�$��8J�q{-R���C�9����Vt"�(��Ժu
���%V�f���� ~呕ws�G��%����/���/�Y�$����^��]u`І�m.���s��!2݀M7�^QIц�A��T_��Ԋ;���?�Ŝ6�2o�]/4�j�@���(E�ԺO�3�������!f}��H�$DV��?prow*�k��7f��J�R�M�^Z�������#,̕�۪�o���RX;W��		~�w �W��G���[��|����̘��a�l�5.��٨3)�O��A9�Ș�=�k�������u����B��RO]^�,;�zUV}���7��|��$c�lw��8���|A`�bU�Rz/�F�Vk�0�T���>W�NŦL�\Z�H�],G��1
Չ8U�X
Y��R��`���޸R�N+.m��T�zG���;��9�?Z�L+BV��t^佐��+ ^����Qk�,0o�C��O�����)ʫ��/6 ����w��Z�6�S��c2�T�I�[Â����䛨b��{�?&�Gw	M�o2�Rp�\�)�c/@ǧCN[�J�<H'ZO㨧���<a�x#������=���t6�
�ci�����b�rE^�\PD������^$�z��~��wS$z��E��,blW]�5? 9�E��`���u� ;S��$B��x�Eu�6~ی���g�0U
�^O� ����%|��+��	*�xO	>���q��$��3�쮣<�r��z����j�Ȟ9t1��W��5f*%g�S!��+�24��y� �Z���*��U��+��Θ�Af��E-t��ٵ[(q ���[�+�4�*[_&[@5}֦�lVP���L!�����Rr��W��g��
/H]�(�5�mO�
ŕ�LcG�pD���L�yz�	�D������Cuj6q�-%�0�UT@+�R�ʦ�r��T�!�pS؞]�j{	9������x8��Y������.�"u�ctX�	/��,�*KER�J^����ˮ]��V�Ɓ��+���΋���$������3.��;�����.ī�H8VQ_��$�DP�<�t����Q���
�Ji_����`ع?e���y����1�Y��@EzH��˪�-ud�-�*/�]F_o���ÔP��t�K��à�qt~ot�1B?7S�c,Ǘ%�ʕ3~�ˤ�bk^��mY�:���R$�0�T2C���_R����cy�R���y��[k���͇�<�����i�0�`�ɠd�fk_��cf�C��![�/�wڧ}� ��vnʎ&9��-�����Q��
�{��˵�z�k�H�kP����>"7�����wb>����;�}�MI��'#g!��$�%;�}������ڝe]�b�IBpC�b�'��߀�C�Qָ��{&������m���͛3�P(���e}��tA?Q�?l�i�2Н��e�=f���a].#�
Y�L��5^��;��?�q�1@`���j�b����M�F8f;L�������)��=t�"1x��OK��o���%����-�Յ��+�U�U"�̐TjzjW�4�
�I^����z�JJk|V(�JG+}bH+�'��	�� ��?��J�U�<��;2?�N��vi2�p�C�Z"%mƽ/��وUv�Q�|���_�P�إ'ekxa�$�΂I�;:F�D��m�_�'"�$d����?�����YP%CC$%b�� &��n��,l����\y�)����H�y�t\o/���E��r@���}i����:^V\�(����K���M� �s,X}=z^�-t�����:d)�E������2ɋ�����R�Z�"��;^o����H�覜�7�2k��LHD�N��qC�o,f"�w�L��3O��4�p�oޔV� 9��%�������e9V:}F=��<�Ob�-�5ju��z����f�U�,�����(�j�W!�h�	�� c�榷񷄈v�;9@�K���5����L�3���X8^5��i��^T�VWr��4O��õ��e;(� �-�T�5��d��B�O�U�B�Z������s�s� �z�/�C'&�ߴ��g�j�r�x%=U\o������I�4=���Q�Rh�C@��uN՘;��͑�7�4Y@�X�"=
������̲`�i��M����/�ӏd�F�v$�h��q�:�=;֎���X0���[z[����՗;��ƎGw���S�9� ݔ��ykVS�S�J��#-������Aɗ���Ltѧ/1W�cY	 �U|��s	�4M�$4��~M侏���)�����]�×֠�Ҽ�x \{/��0>�6۴�x��Q> �W�K:B�l���.���"���Ι�ʠ�RN3�QP��a�ؔ�}�j�+���s �ڍ�����)��=�W<t�x�-�8���t!��N�?�ŚE>���r��Rf��O�RE�%Գ��ih�{&�.ժ���f%D�䔇�f݀z��ٓӜ�5�=�����B��9qb�ucj��&�-��Q���"*�X���/��iu�h�_�O�/0��eS��quh�bz���o�a���x�����j�1�$������&Kw�[٧�������ل|� �=`7JV�����W���H_��r�~u��J��|v>{~���΃�B����O*�����]# �C���V��B�w�s�"z���N8m�Ű��º+Y+����F��JM��TϽע,��gz硽���E����쒝~X^��Z
�t�Z�������X�G�بv�J��Jjj�x��rlW<W��)�P��������Q�_�(~]�V��M�A<���T�L���|#�yH�>��G�8zQ�ݪT
��BZt38�=h�s����k��`
��@59R�Dsބ�&�9���I�Ȃ�����5����������/Yr]�%�ԫ�ޅ���K4���ÒS�?�WH�1��z���7X%�_�$s/�oպ�q�u<�
&�p^#��F^��= �.h���P�_���?/�o6�{% Sp�7�w��硃b��y^��K�
X)����f0۵~�zN�!16|} S���7���{>�����R�&���'U)�uX��%�TRqV��C��1^�/�y딓w��sZ�N�Y�@��T&0aQG��j�TL�����h<f9�p���ˀ�K(���h�����'��d��)��`\r-�۝ր�Ĵ��M��G�w�<l��?׫|
���xQx��puv�d��c�)l&�q�$�h�
t^�(��_�H��kxg��y�@�����"�;\�c����1����;!C�!�	~O�а&tz���h� o��l���)���:e^��FL{T2�Sh��8q���..K=c�"���J�u�:��)�L&y�����y�+���W�cC�p����s�f@��]��J�俞ь(�d�_���>�p�K(p�7#��uRX��-h���^_��"R�1�d�:��V�����k��( �#��[[�ѕ�X�b��yK{�L?o���1F(����u$�^^}��� /����mPPJ1E
N$�uď�>3!27?y�)i?���� �~��-�}c��@�$�u�a�b٧�CT�T��{~H3]
r;�GM�Y,N�yf��'�:��%=�km�"��;�7%�9`�B6Y3���,������-�.��>F��E� G���ɇ%R�ű��H���p}_��utu3�}��wET�r��LL�x��zȦ��������d���|6������.d��T-�2�5�-����s"��jp��ݻ�u�����$��}��)p���XM�Oj��υ)�U�J �����cx!qFx�p�w� U�W��f��<���[�U"{}�y9Ylf�>qX
(����䤎���n��e/���zk�s�!%�` �R����o�~���l�SǢ9ƣHf�O��w�9t�ֵ�����	܉�	8���邍$b��.[�]�w]���4B�6�#�\��ZKOBe*���!��/vlߌF���/:�J�LGF����w6�C6��B�_�,^���FIb.����(���_��o�Qh�!0)��Х�ߖl2�#��-k�$�<�4���r�ՀE���?�?YҲSc�E�ʗ�+(fj:e����-^^�����Т�H|%�\WT���� �0��4�q�q�쯴9�HS*Qb��c�Դ��Dy
Xk/zƄ:��������g�Պ5D{n��=i�����p���,q�8;%w=�G_���ש����(i�jkkK"4>6���]Z���W�`P��kA��<s�M��Rfd|5�'8	�0z�!A�SF�염S�z��P ?��T�\��������Sh���a=������U�4�����ݦ��B���;\�R���T��c�����KP9�T�	ȇ����Z�q�����^�p_z��� ��P+�m���xq~h!�fd��v����	9yK-�������g:�Lo�
=�֮%�P��e�+C�R��<��e��{"3��03mw��j�1:Ҵ/��]j�����B�)�p��!���9�y�]�r�{m��n޳)��e`������^M4b�ob�Ѷ!�V�S\�}�n(��F}^�C�yU���;���������׏cZ��ʾ���c�P�<��{<1�G|��λ��26n��;Y�{�.�S縼n+�V�3��ж��z�Y��&�X
T�ɧ�Es�G}����U����(R�����1��V?�� "By�סױ�Z�8���(�c�*4��i~a��C�%:�߿� ��6���._� ���2����dH	u|B��ǲ��,�����;X�猴�m�3�YS�\���-l;B~AaK�<�^��V�
��Pű%E4�c�t�k����Z����=?D�W��j�:#� �0��d�c��бl��5g]\�~܍���׏��a�n���؜i���VU��L֍j5`���w-�s|׼lQ�Rm]u���7\�>~�u۷%�����h`�L/}�.umǽK>�掖��l�2���wY�%�-��j~��F�zJ��9��0H��=O[�,�<pV�m�$�4A�?�s�p����Mx-ٮ�,4㉉���>�.�7u��qu������������ SdR����f<��3�,z联d���'�Շ����0秀��ׁ�'�),���s����E���`8�O�h��+��-���.�2����/W�O����O�d¾,xU��:e��X����謃��0^(Rܵ��@(R�=��V\+�
ťX܂K�/�"Z��;w(��~d2���{����7g�>/ǎ3�^�R�%|�Y\|���Ml��
�
�*nd�v���m�VJ�$nb�+e�@s�L�W���So)���P�%55��B�6f�#�ַ��z\�ͧ�?�w���ۯ	I�, Ptđ{�T�kB��k{��	�0_���Q�Z�0b����%=a���Ē凉�#:�7��V���Ǒ{�m�i㻵�l���|D�%<��U��>K�͵��kg|�~l3��9y
���]�L�J��^���_zkv�$6X�.e돗VɄ���*�yc�P��?��t����own�d�N���;��PĪC!+SAQ0��z��|�
�sP��D���f��J�!RP@$a����N�`4ʴ�튍�t��ՊBW�9[I���!n`ii=���D����K��{��x���_//kՏ�s�E>dĔ�g���Gڧ3��Y	6�cW$C[� r�C�cLU[�����4�'�F����ΧCCC�AH�g��Cr�����)'��.�_�h�	<@z�D���2��7n��K��ESD�Y&��J>\v��^<WǵB[����$�B�7����z|�S��Z�{�s�+ ��^��M�9���T����C.I���J޸ڇ �_r��(�$�C���h�i�Һ�}���� 	���$ 3!��X�<��L����p!J��1X��������)�a�!$]�h���vƹ�V�ý�4�W��`���E41.{i�<�]:4��ޙA���Y��7Y3�q�瓙U"�4��W�,�����.�~&�&M8]�F�LZ_/�����@'P������=������A)�i�z�{��˟r��0J�>\��JP/ J�ih�ʑ�]AEss���"�݅�ʭ�=YgI`|]\�}�\6}��;�2�l��E9L�s�h�;�6��h�>�����&�A�܏����$�>��l=>�]d�;tl���[l��C���B�t
��@^��X�%��)V����L�0l�������U��w"��������4���v�Ū5%1Eq�8�7�������_�=�w̏E����,�NA~,��D6n6ٿLq�j��f��~����ߓ+<������c�H�7��$$��E~w#Ltb:5���8�٬z�pf�	���y0E̩U0��BǍ�U�#�]e�)| �����7����}�)�g��L��#vI�g�X���$r� '>�P!�"<���<C�2-�6����T�as������r�N��i: *k��?a@T�o�Y�+�e�Ȭ�ގ8�����H`F�� hpLM���j�=k�wR���l�(��� ׍��6GP�v���EiI�9W����X���1��ri��o���Qkγ(~��[�K�����T�T��M���Fw�M~�nY�5	�^9��h�b[օ��E禵u��c�mW�m�A·���$U'�*L�������V�ąԝa�eQ[Pb1�����+ �ܝ[��7��J�M`\k{����̥��ݕ�dI��_���ޓucn��it��W<��R�Xǝ��_���Z��ݬ:�:���9�aD���+���UT:���*�%%�JrW?~7��P*���V7��M��:wk��sb��v��YZ�<�gI &7��K�J�3  +q�|�����\H8ܒ|\�^(����i �v�`��7�	�
B�}�i^(��~B)ߣO�G$�2�F���ru)�\�߻k�YrX�Y�9}����������b9��Y��|�[*��Lu��
H��B{���1��)+5����B�Ҽ^��q����.<6��O����~Ƕ�����XA:�� �%�E礭f�!���< {IZ�bZ��/�<��Ko��̠���#�o���ʫ�a�P]cc�Ei�ڰ�S��0+��#4�>n@�w����H~�q9ww�66���,PFňgp)��'�!:~�k<�:;c9ϲ����"?pQ���W嬅�.)'��mj�}���-���?�r���_!S��W��#��_����E��%LӻO�?g�ۯE��x�mO8�K�A�XsRgj�~w��t�`��Q%w`s����)0�%~�5�S~��3i˩Jj���-�i2���6������w��+ďK��w�j�������9s�o�@�x���}.���gf���H�K�Dh�pUp�ACh��O�iɗeC{4��K�v�F�T�8|�\��=�@n��A�Q���(��M�N���88��O��[�Z�-h���M�蔳R�F�x-5���8�VE��N��h�E�Y?&Orי�1��C�b���\Ɓl ��s{3	����d�6���u�b4ol���Jv��Ti�-�w��}���{~ǎ<ӛ��k��-K�5��`=�H�qlr�Sce�t�i����`��`��
(C�$��U�&�#�"�onn���N�00�շ��6.�Ne�jŅᦻh��k҇ۼL?]?J���� ���������Hh�BDkk�+-"e�ɿ&~��YF�Ñ�XќB\k(X��E[JC���1l��m�����B7�Q�ͱ)?^m�5�b7�s>�8��o:��;�na5���M�O����|Ӈ��Z�����tT�tba�������6I�3�0��R��T#x����)�&Q�J>����ޙ������JAG��k�1�+CQ���Q�K���2dv<���˿��Yߌ�b�����*�ǡL��C445�Q�ا���߄bxS�O�U��w6ƈ�	W�d~d��j��D��fl��s�җV�&�ԋo<8�bJ��8���y��t̋,�q4.V��x-���/�=�,[�o^<�;�Jj���є	7sZ�I�\+����0m�4��RD'홧�]�ͷś���?z���=	����e��("�YQ���_�kʤ��Mn� ]Z-�4;K�ӿ(�r?��g�U����x�)rn����+�4����%�!�/���������z_Hz� �}�\��{g�S���;���+"�>k�؅n�S���6�{G����8�_c�^�s�^ڢa���"��ܼ# ����s
0r��r��$L��f�Ε�Yd���
*��59H�&���W�t�/f������x�^���.���g��q�M=�]b����ec�������~����E�W���^һ	�2
�85�M+r3��du���Z��]\~9*���e"�%�ꈞK#5�өt���V��pFw��#tl4	��=!�ψW�w��W1F���w�=y���l�k�CPF�H�tk��:ܒ��W��{-�f'kGg�7sJ�p�{�'�j��V%�{�kC�?E�i�-_5�aA�l>���	ףQ��#,#����4���3�Kz��I<;e�1@'���K�%�EK/����o��=���Y>��	T'ޥ��S<����U�OnH�&OO<zK�ua���)��2Qb�X�%0���w���/�Is��3?]�z� }\llъO���NZ�w̕���AOYiή�@�~����MP�b��������d/se(�� ��t5A�F�������E'�TJ9Fٚ2"g�M��2�p��#��O�.7����u�9��'��� PA�W�V@��n�
RJ`v=p��톀RZq�B�D^���_�疶�=.D5��
���o~���R�&��j�g>W(�6I(�ׯ�����8\|}�ښ�q�Z������7�S��7�H�/ÇAC\2t��'x>��a��'x��t27�����S⇳��ݬn���ݩ���ߍMwsm��m�b����_�,�ڸ.p�K�Ӭ�����G�-���>��l\ν\
��y���.������a��
�!�=;�B�w�;�L`���ۋ�*��J�� ��np;:��(�iqO�R�ځ4��1�k�����u`F�r�N�]I�3�G�6��*"��\��C~X��Q_"�У�{+Xζ݌[S�cQ	���� ��n�i)��2�G�jڳ#�{~L����.�#���<��������lȓ\���dcB�/X�d��F/��}ɯ���%x5�~
����Y�F0M/S��揎��t��)?��mW:�z����<�J�/a�U����jwVM�B�jޢ��n	K�6�c%)��$���I?@�۞U��]Q._���ȶ�`I�޹�ujR~!/O�l1U:D��о^- �"��:q�e���p�M]'*�<L��1F)Q�qp�%8&��7�k`j�$����MF���,9u�����%Me-[��s�h�u���Gq=���O�.��f���S��){�/�ڜH�=F��Q+Afv݈��X����6鎀T�Q�o�|�����r?^ ����JY���# �u����5ii���*R�D�::_�_��k6y�	9NΫ����xw���z������ܬg%[k}q\; 6T?>Y�E��������b���<�tN�� ����_H��ԸVP=�GZ�Џ:7���;�[�O����ρ.�G\~D��M?0(վ J��PB�����,����KC��Ԕ0R���[i�u>2]��,�_�,��ρh�����/Z(> ������\�j0`�揵����+V���!Nc���K#�g� ��I�.	�I&X<\�³�_��_���-�;
��?02ib�&�RA���E@3�2x��$;|aO��[�<Ѯ�S*����/j�V��'���̥:.)w2����U\-���+�+�nL��K���/�"���j_�H��?�f��pUYO↸��c*�����H8�vN݅Qޖ'����
%�.�0�����d��(��Zo�%.���Rյ"Ub3I7�t8�p�]7��N�X���{���.��	��	�Hv-���<��l�lft?d��������F��S�cY����@]����'�,O�����Z�F:�a4�G���Ϋ���T�y���	�Hd���==��H���%{NՎ/D\<�TQ�o�'9X���9|�+!��4cI�%Č�"��ӱ���ζ��d��š�$+7W8�7@�B9�.��S�5E]�ǣ��L�[ہ�����k�,��Z7B+�X���x��v]���}�r��ȯ�ͅK;�T�Nl��|��Z҄�*r���_zκ��|�`	��b�H��5����rp�U,���U���<���|��B����&��:K��!&��}��>Y/u�k[OlR�@F����(\r��5��Ϟ4Ar�{�gv�M�'wr����	�)�l���|��.��� �7� �b�:�'��W�����9Sf��~ܼ��Bc��r���U�(�j$L[�Wvl$�s��_ܬ`���u�Q�t`#c���F_��HU����T�� ���R'w�D
&�A�+G��G���U�Bz+G�z�.|V�e�Ǟ���S����s�
+a�E84�M��Z�+�����8�'|g�g:T�c\A!�߀�x�$�0=���y����a��j���@����,�ŝ����M0{��Jx�0�G�X���L�?�0�]\�����&�x7G>�j��~�:���gKo�H����w������T赤CK���*l`i��n�p�oC��P��+	���VMa�}���ɈQ���%��;� ��OoS�P�2ƒ�B��u�$���e.�JG�rȴ�g3����-��|��������bQ�\|�B-�e���J��*�y���C�5 ���+ss�p��� �����w�6��n���Ue�+�"A\Jj}�=2�>��3��t���oƜ��$}xkw$��"���@��,�ڙJ@n�����M+.*Mr���SV��񞞛{䯣�Q���ک����;�XV1@&z&66�yC�UT����Km��}66���	=�Z�I��y�FA7r-:���͖�:&0�P�,~��FR4�(q�<�3 ����]��Oo���X#(�����X���
|�}�>n������G��~w�D�J���S|e��#��~�4X�_<{��"����F��s�Ю%�	��7 ����/۬e`���X�y7(; (�|���.��=�:�{�l���g��[��z���GC�.����X�B+4x:ɱ�mB�v>#���Z(in�7k[�lEnϞ��4��ӤX#>��B��*���)pH�k�W��o�+
�gڞ�˻�j�g�k8���p�)\���Z(C�>��j�L*�aܣ\��>c���#�~�\l����va��xr�����3�o6]0���g�u<4�Wk1���b�_�Ys��`���c#��g��0�2�ڨZDeʹT	�2���cⱣ�{�yDJ�'\��O�ϙ��Ϳh����y��ƥ��}S1�	vU���X0��=xφ}��c�4}ا���?w��/�p~3�qi����ށ��4��ׁu=up>�4����|��g�ŏ��r���U�c���������lbII�*�֮ߦ�MAk877{{{#΍`��I�&�®�{!(7s���b���$�b�W��Gr��vq}��W������lra����DG\R��7�㳣����D�9z(�Tº��^A��	�_�@}�@p��ʔ��JƘ�E]W:&�\m��s�"+ڒ��*�#�4W	�?�R:´���޸�@o��B��I>�l�oTV��ƒg��D^�2���r�N��#��4G�*"-��k�:PlUWEu�Q@ْ��1�����R�̄���ے	�.�8z�}��&���)[��ѬF�D�*먪����n�3��𵆓��%h�	��$�[c��g�i�f�����ʅ��f@7��[!<ں鶎q�&����L�dE7p,�+�0xf*D)R�]��iؒ�#�y����?N�B����y�R�m?T��~HP�n!�Ȧ��,A�o�6��09z�m�����:Hy���Ys�����+�w�b`x�?+�֢��|w������F>�z�!_�.D�����b�7��Y�?�n����1a1,��g��)�:Ű.@,�n�o��MJ����h��*�c��W�{a��7���Vyl�z����B���~��c�/���^�1|�w�SU�[�f���N+��L�Jy"?@�0�8gs8@Ue��5Qa��n������*Gj�_�l%����g�8��Uⷙ�;Qv��!<�j���'c�v'ن����O/R:���M�w�UL�;pqeee=3zp�=�ǋ�	EBG^���^�5�b�a�Sd7B�Md��^�G��T�ƭ��O�s�������e��Bػ����a�Z"�^b[l�:K ɛ~�'&�z8�ZY�:�i�K �!�ݎ�c�Y��&�e��ۤ��CԶ�U�NT'\#��թ���]�JgLZ$@ʉjx4����.jꧬ�%^�+532لObQv�e��f+L<B��q���7����	�VQ	~Y��|�тgi�H���r�;=!}5�3��R��\I��ou���L������1#�����w6�fw��{(D)g~�T� �s�i��0��?:���KJ[2,m��l [�_��ABc��8 즥�ǖP��w����N/��Ul�������gڼ�Zi��+v�8w��/�6�н}7�s���2����-�5�S��<��-�_������E&�t	}q�\�����K�TLGR6i����u��ru���W��̊�b�O�%�eq�%F6����M���Ѩ��Ġ֧��Y�=��1Pc+r���5}���!�q#Q����hD��ED��v���^��5�*v�og�5����Wk�a=�j�ն6e���Sۿ���7��-��.g7��v/'��$U�����<ћ����kr{;;;�Xޡ�}43���u����c�t_�[7	fk?b]ф3���.�w!�1Sʁ���w�`T����J��D/"ˈ2pyM/���ǌ�G������l�]��C{Wޘ����T��X����[�M,�(���'!mv�)V1��O��V�����1b�n
=0��@h�>+�����EYE2����#���,;3�'��m9����!ѭL�+�B38 `v'��u��Ĭ�yEEE����:ӟ=�����U��z����R��9J4r@�Mw{�ױ]6�:������g���>�_��]�~q���.X3O�j !1]l�>��5��n%v◮�;���M�ӝ���2�.�\ߠA<�{i��M�7^$�"�ws�<���

����Sj�2���6�a#��?���
'���,�����֧�w�j���zxg>�n^}f:��]ʛ��Y�IE�w­��3��N˱����@m�����ߖ͵ܻ������#��~�c���t�@�ɱ���dL�Ad�l�z����s��.t�a�юU8�_g�#e��2�R�;Gǒ���5l{͞���g&�3��س�$}:�j(&��x�vӎ�o{��ιz����RXɵ����X�suS[Z�D��`��#����������n@����S#=� �QNVd/�����<�*��C/�fg��;�sM�$��=��)��[�tkg�H VS��7zM������c�*�crBt�4���\��Um^{�qX%]�UKL�[v$)c>q)�`��G��~�����p��)a�e�O��K��ц��<y]�~���N��c��"a�^���%�=�Y���;ƚ��+7��?95��d���2�ݢ<K���{���uH��e���D|�?��=E�K)��]Ʃ��z'��7��a4$E���zD��F��}'�.��Z��갿�a���r�n�|�����>��L2dH��Ty��p�z#���7��6�mt1F�MU����#)��FQy�m��u�k�˾�v3*9���{"!���jL9\J��ŀ�5VA��I�	��늍����ޣ�4����c#oѺ��U�^�˅Z���iv�9�����#!&���Jr��x������{������s�P� ���[}���2�������g�v3�w�We0V�tϓtk�V�G�a_ǰ�?����I-J_=o��O^X;(���QQ�^4{�R��|�zg�Y>#S�,�6#�H��z(��7iw:R	��#�S-)�zc�=@���`(��/,�o(��[�P�w �_j�o�R�g���E�a����%c$CL��.	�SX�Rr5z㯣.��ұ��a���?�A�|�ï���1���G�Gڀ�m�b���Xk�O߰�n�G�@�>Eh���k�VD�����(��T}i���,�%c-q4\�i^���t�dSO�𥒜�p�g�O �z�j�މ~^"��S�����1?v�ZI"⭉$����6��{���#�K%�1�6�1��`���T�U,:п٤�lH�9�p@������?)7�ŀ�5���3��H�y�>p>	i��tY��XR�+J,ʟ%�WV�#�#Lq��l+�P���cV&?!�-�J8�&Ҥh8JU�E��*��7+;�fG0�«�������k�Cc�Hoݳٳ9>�7�`���:�2N�h��9���P��֌+��'�*��9���ɿ<̢�R���O2yK�2��"Ήʟ�#�#�)U/7�t�c��Uࣝ��-u����3�)	�!�~������h[0w2���"Ak���w�;ь�8�5�6f�(��Q���p�.���P�8p���2:x��_���]�m�{	�>��N��������K�pփ��֍��z4^M�������%�,���&����=��6���ml�1�b0;
�;+i�x�[��M�яET4~3w ���4v�Y7yo|zۨR2e��Hk�R��� �XP�����V�2����w���O޸2�{|JWt|�#;p��������w�^	|�w�e	И��ӍX]�9��Wl�3oR�r���Ŕڅ�%�ұ�s�J��o����h����~z��x�
ˆ&^�2��
�E���>j�酹��
���9kYGcV�-Q�_Z��[�V,����#���f��� ���+��:��f�Z��D����.%\���dVD����@^�?�/"
?�<�}s�_����:�(��v�]��m����4&���P����l��j��WJ'�W�B�lrq����7��Ԝ9
q���LƝ|��㔚ٛ��~z�3ޙ���5��8d��3����S�u�%~*DO�������VGyŃ���dz����?T|Y.?�7��3α9!$���T��^��M��j۠l_Xf���@����*�N���!��p��g<���ǿnSV"4���d��q'�&Y�p;��Y�w�l��{%�H<[�M4]��m媋o��XuWxt�',�W�ڗ�J:�7�O����%�͇�B�a��74I�xj�ɰ�v.jå�r"��bі�0U� c~��C��O��ﮏ�sq/F�#
#8��yԴG�=tpe�B��*X�r��ON����]��9Xk�U���M{���jn�|���h#=P?dhG�yeU�2�O�����l�+9�?5��v*Dv���f Chr"�䠚`َ�|xc�y���

��㌶���h5K6���>t@lbGFR�Ͽ偨���k��%��}��yo�����i��_:&���rk�.���z��e�G�T'�{T~5��|���}�+�yvƀ*��V��	rp�_�x �}C��[ݙ�r�ǰ�B���`���#t���ҳ��H`�*i��	���*�W�Xp��쫠�2�Ǡe�2��9 ������/��<JB�'{�h��K��!�7ia�D�c����;�3O���$]L�0]������Sq	���X4i�>ӏ�gN����է������RtJ���*����EZ%�װ��~�=� �O�R��f��쪂�E�1c{bZL �o(Ɏ5�%����W��[ 9����.��ք����ds��	2QD���}�:8A���r�E��[	������1ZkRfM*�֕4� ${8�q�=l���}-a��w�P4�+�B�*s_��z~��̠͟ �qB�4C��Y'��al�UD�T@�I�:�s�L;�]n�";��kPjvЎb�Ŀ�Gt���k=�:����f�?�Ǖ%S��:��p�t<\���{�|��ӗ��(�s���0Q�$T�n2�N��_�� |Z��~n�e����Z��g��y*;zx����`ʧ:P�M�BX���rz�ş��o���L���֚R���N?��|o�]�a�]��-��'Xt[�<y�>�p���:=�xdʴ���������i�U&�ۗ+g��v�ɶք��AP�a�CB/g���MT�j��RRB6L�D{B�=ڇe��HC��/1V3�\-ԍ����>�1z,��X���(�}9� ��̓�rr��
x%)��3^���8�	zy��Q�л������8M�$��G�{�mk���e��m�ܟ���e�𱤴�6��x�u�tXq����d�*�}~��x_��v�>���?k��­"xg�*�|M��U�lv�/!���+Ô-�E\����$��*��1���0�A�=WyZ��+�#ĭ���<�G�R��a��j0e��/��3O�HH���t�Gr)�R�4EZ�԰!
n�fHfZ4��x���3};�� �*��&� Pk�/>�LǛ�"%��#ϖ����b[Sn$q�3!y���
|Jv�%?�^|�Q�X\&��w�o��Ԑ18��nK�/���W�����4��T��&���gz���9��� �7I�uA[�G�γ�3=�=�ܢ;��+�F���:r07wuр�ޓ�:Q:�.�g�?판N�P�m(i���&�T3�d��3`�����/��E�di��=?������M�:xd��g[�~4v���O��nд�Zt�}��KUU����K�g���$x|QI`��*H�����Y��߄�8o�^3.1y����q��a�~��^�6lH<|H�C+�=����a]��7F?y�AӶ� ΃8�J�;���qW����cx���x�������_���Sj�'�ȗ�kl ��C��J�%�+5
�����a�������;��0�����z��ҿ2*T��N�r�嗈�xZ�]������Ό�̹o2O'X�J��ƌ�6Nyo?�R��*��P��|��ש诡u�g���x�8m�pi�`+WO�/����e����	@�
� l��-I��~/��Ɯ@e��7�H��a��݀��ؐR��k/��}�����G�L������q��3P��MF���O��L�(fv�ns<��w��O`�|z����֪>��;�V�mjU�����H�t�w% R�?��3a��paÒ3������@ϳ�x;� 3w�]v,�{���%j@��V�5׸�R5U��D�9q�$�=�ّ��f���V��/���%3����/��
��J���n���3U�[���ִ��LGKa��*LV�=h���P�]�y�3!��'=2�H#��z�btv�d�$�pp���%/g:&7�౗��쑃�ݾ�qz&��CA��!�|a���>�cew�	�,�	����	]}�8���H�������Pj4л���^��,,z�]���7C!��A��'�v:{��Z���	�
jp��'��p��`s��#��3Nn�=�n�����L�9[[e�����4�����6�a���6��t��S�,�E�� ����7������?3��a�;�x�0�r�U8C�!�e^4bDa���t��7�'��*�}�X?��mg-]_�L���	��@��o��.z��������7�d��J�J�s=�9�}C�?V����c��[�#��~�G�R��I����n�՛��~[/b�V�Fﷆ^p��*UY4w�wbLU��-���N�V܂�(���5��x��k6j�	��N�B@���}�3�䀏���9����V�$f;M޸��m���ۃ�Z�������e�+P�)V;�����#�<�9�7Z���Rl3]X���<��,�����f�-~�qI���sˇs,GP�Tm�ۖ��+�8�ΙM�Lu@���z]P|�O'��������僋tG@��*����%���P�c
)���+)��[��e��籙 �����UN��������r.јtxB�O�w\�voB{֓Y_>��}��L�(秐g��5K��P�)��Ey����)��h2��,x[�Z_$�Z��S�^	sb�����*Wh린S�Z�І���U�X|I߹��,��vA΄�pĲr=�&A����� ��{ń3ji�oF˗0�;���ʶq_�˕�eL��d�.S�����j�o2���%�@V�o_��ݑ?�.�3�U3M��ir�Iz��ϑ��9JV��,��I���D��T���$L�}�����������U�g��^���s��#��l'�Z���$v:Z���A�̯��(r�vJ�t�h���оd����⫊���^MJ�������>P�h
ŗ_0;��0�X�`/�y�|��K���7#R8k���`�����\A���rdp}9�켰D}k�ر��<j����oo���H�>M��,��z^C^C3�1$'�� ��X8SGp ����?v#�������S����q��!!��\�JF���O�%Q�I(�S��J�:�q'��6s�����΁ˡ�`�Krhq�/lH�PRr�B�VRή؜%��9w�cJ�v:��S���YX	7s���ws�m�vo�ܛǚ��Y��������W~�eZ��vE�9�~ VJ�G;�A������� 0��,���}L��7�uvb����`�WZ75��!���l7oeɽ�������3F�����7"-is����6W���on�Аv���\���ɴl~�����<�����)�Di�}PKU�`�t��U��#�[��H�]��1=!�UuH��l@!q��o�Ҽ�����s����J����Ͳ�FB渋>�����c,���wbS�^8O[
������+�W�~vG2Z��J�,��<�Cd�)1=ˬ@�='<�n)��Y���(��"�.��i<���~����F`����2��̂�G®���ŸU���?j���;�m��/
�(��A�ߨ�>�ٙV�Y4����ra6�ۯ������"h�k�f7�	(��Gm�^�M"�"N�-�������.`�5�?��?6�)qX>f�Y<��J��y�wY� 0$
���%?sKɅo�Oz�'[cm��-p��.���ϘP��4����b���z�ڃ"��X��$bA:��}Y̴s���[��с@�؋(�grR���o�G����_��:s�A���hml�uJ����<4c���U�V������A��F�<�4Z�Q��!��k-8b+2o�c����y�1kHѽ�!�.�VN�bHQ��E�ｖ.K�n��r'��-ԋ�|���~��'c���5ͯ���5��5m�j�)���FҤF{� ����@���`]�v�B�FC�����h�l�?0%��� =i�q�-͉����Ӽ��5�h����.��5y�]����F���Ř�J�+�Y��%�����������J�T���*!g%���޹a5В���oq(>-z���	����k�h�ѿ�ո��b���/���9>��Sn�jPZW:j���tl��4%s��^+b8�~�ύX^Pq�������]A�Bj���2��b��6&�;��sPB���R7��|-���B��LW�������%6�Ypp��K??0V]'�$�G�A� ����D�t�å	hf���k��"���������9�+k/>�h��/����Ưy��	9Xu\�&`������a|q�dԇ�Ž`�C�vwL�B�1_?3��� ,g���\vo����i�#��WW�89nS�|X��U���5�A��nA����0�������|�ȟB�R㶶������N��~�j��:�6���ϧQ�w<r�C���LP4\��)���PQ��m��'f����ox�����L��������E�|�z
��vP�:�dO����t��y�l~ԙ/����j{ʘ��'��$@�hƯBgi>7���v���D3�*�<��l����g�*��O����+7�;Z%D[;���'�W!��AR�'ju��Y��	_���c�o���[f����z�JG����鹠S!�89������U��2�8n,���"#�v0�9'?4�9�"����}�����%0��-q{�6㚎MQx2T )�Yv����9�UX@9)��fޕ1����t��M��"k)���juf ?���+_�����M��9��Ɛ���h�b����V?�}]�}��
۰L�_�,�o��ս��:��ʲ���<��Y:����������D̀bQϿg [�k�ћέ��	'�u��R�O�GH8
�ڕfw��p/K����ӛ���^�i���4��Ƥ�5�J�n���,䆡�>�m����~r��-���QbW)��� +��z�o��o�7����3�UN�B�y-XCC*���+@bޭy2�u��>�2�ӳG�gi�JtC�m���8V��G^kJhfn���ϰ\��x���E�D��;�����L����rx��^�Ja���"�q��Fl�D�ZU�K�,�W*_]��l�����{B!�zS'���l��y��|�V�G����=9��m*�Z*T,kk(��ü��e�ƭ�n�T�BՂ���A��Ɩr��=;믫��'�a�3r�uoR��Ja	o	��t[
Ӕ�X��d�U��i� _x���%���j_ڌq ����S�"Zi �]�y��7�KH��R�]16:$��@].Τ<��C7�}��u�������*4�@�75B�O��0��<_!�[�煘�w�,��hQY�:�K[���'�`Mqі��-�Q��7����Zݾ��M����F�������(�f���@h��jF+�� r��5'���O�������5��8��r�����;	Wk��4|�����<����TT]C�(�J)�P��/{�;Tg��R��r 7�V�C�TyL����R�7�3/u<���@���6r:��0I�P���]K������`��w*q���7z�pf�>���I�J|Ð�',�g�ϴHp@�S�B�\�A֬<�Tp�bfff��T�o���|����ӷ-C�b���욭A�`CF-±C*g����t:�oT{F\�@�`���0YM%���I�Z�]Қ^���yZg.ŕ1|�ۼ��u�X��A�W�b���c��t�ޙ�y��&���a %q�l���n�N�9�P�󫄊�e�";��Kըf%��B��~��!�����3@ݛ�Ș�=%-HG�X�T����@!�S�8:�(��Q� ���M�yM+D��΋����x��:!HQ��Rpc�ԇ()hY�j��\c�1�Wc�e��!9u�$"�>!���ш�浠l�p4-|���A��x�y��;_9�F���	���Z�h�2Ah*��v�NiA@�A��BP��#o���ė�\V|����ѿ�	�������?�l\r2�9�.9�xNƎ�I�����󊣳R����i�d�8������s��y���q6��3��4r:��M#G����O�<=Yq>q�N�~~̏����������S�=8b��ko�Eᶋd��8�T�y1^p]$Y1ћ�"3�k.�MH;֘���d��VLl��K�1�ޘ�zâ���*�T�&\��H$�����ܹs�?���Gw>�;������Sb�6(�0�X�*5h�Af�1��$wCd{k���}�\�ΰ�C��\��K��tz�����;��q��>��g|����NOO	ё)Qڊ�X�N����Z�u
}_H�#rN �<_�J)R�2Z�r��5nܸ�����5e�"xYִ�-�F���_�����_=��m���1��F���B��R*�oX�J�F�J�Se���Pa
�|�(Ć�G���HϠx�����s�T𔿂��g)1�wm��*56)�@i�mR(/Id*4���&���4!�xc0x��uN��
��^|C/�2iiW^°hɁem"�
.�wҪ���!zB�00FA�r��zŗ�"hO�Z��W�����>�����>��ޠ�@�eW�^ZO0Rp$���оК�+��7"�yŽ�O���]>��]O�9[z&�d��,���4r�Ԍ7��Rs>��M3��ٲ`��9_h�����|�s>��5糜�a�0<9�9:��"c�4�ι������G���x�j�X�U&^������b����)J@ĚNܙJ�t�b�����hB���(��	A�Pt��`�{���Do�6�����������p��q��}>��9�~�9�gǸ�����6��2�ŋ���8����R��v����ۣ�t�֧���*�9GGGܻw�����?~̣G�y���l&�U��))h ��� 5�A���z	%�{��y�.Z?��f���W�0�
~g���ϒ�xJ�\��V���vi�9�-�S5Ƚ5�A��eNx�zC�@�E6�%4�bs�!�N�^�6�q����b��|����;@�
��_Q�H���HX2�u��i-mGA6{ҵ~����_I��G��^�j��*U�@cJ�O�GLy���Z�-���� ���"uDWK�ՄJ(�H�2:y�͹�|H*1X���:�S��i����cʇF'�N�%列�"'3�?	G+8bN�7����g>/�L��5�R�ūl���9�T�% �LcQ��2G��g
0����#� �(A�c��t�VƳ�������l���$�q��o�X�RU�S��"�M��$r�I�aY&��'�����'l�	a%�g�������<UU�X��k�b2]�M����^ �*�F�ֵ�ȇ ���EG��de0:E�Y*'��!Ja��j	��EN�ۦ�jc�X���2YwR$T ��b��t%�s��S��kD��=�Z��sr]���Ŋr� ���I\�b�(���(��r���Q���0Q��>�ՙ�H��ڹ ��f3>y�ݻ����>㳻w���g<>|�t:�\Ք��%&��%'&�T	�U����/?I�#-�\[Ϲ&��������zE	���!U>n��ͥH�/$k%}�s�'xV��_������H�i��u.��ނxoZH����:��Q�sq^/�=)�>�P�)�r���R#J}]�`ĸ�7�1�Q�N��u��T��&��u-��A{b4��8����Pr�^pY���M����:��ʤS�S���TuEU	L_�*u%(GM42o� D�,/�� ��{&zq��rs������H�e���AA4�` h�Ω�E�J�ƩH��V�ZI?���Q�����-�!�sr��mMar�N=o	Ci-�x�JeT��6����dK^<|ΰPbyE%��J����Y�Z#ˤ`3��I,]L��@+���EG��ܿ��'j'��(BU�5X���wiw���]ZE�"o��0d��'���u���_�h�v�	�:�\,�+'�M�ʳ�+ `�"�RA�8GD�Ȕ!7���[9.�dQ�Z�5UB�Q�oJ%�r��Udt�]:�y��a�
���ڌv�C��#�lb�P�բ�s�JFM��A뒪\0����qrr�����x���)�ɹP��F��[�R��F�����#���y##*i�V\�rR���/c�x�b���4�m\8�"����F�/��o��_=d�h~�x�>A�m�|3�}���q�x\z������4^=��sb�V_;��xw1���9ɏ:�{���ʍﯨ|-Ǒ� �'��U�/S��������k�>G��_8�B<�|�G�v:Ѣy/���iB�	A_��y�<ޗ�J'����_̭�q/��Z��~���s���'�`2��	���yKP9A*,C�2���E�����h�KM�R�'�!M�E-�|I�0e3t��$�T�6}�Z�5�ב���uE�iUR����R(�V����r��^�l�r�b!�W�Ś�n� �Rh#��ro|�y��t)�V�r����[�G�����C��>�^k3��"�Ԧ�CyMnE�e{�M��'�2��(��ȳ	@z13ݰ����v�`�3��գ���m��m��v{dF�!�L�6B����nwuFo���hk�<kA�8/�,1]S���i��v����t�V���,ím�v��/ݲ�R#S]2�VLg��e�d��QW�fLi H$6��� �m�o�Ռ��˥Y\r��K뉫>z� �,)W� �k����ˍ�˲d�,�ʊ���~i��86^������x����(� p�dH֍��_R�2�x���6�И�; �;d��Q��c�B��x�h��Ժ�&h���JA
g�x9��E��e��W#�5�	h�r�w���h�S���h�PR;L4�R�����cNS�����b>{L*���z��?���v�\�~��7�bw{��( ��:@0�3�^H��T��0���fa�G�6�0�G�W7�����'O�p��	�{�K8�������jv���r���P���܈���]���u�����sNON��q~.@�/g����X^?�0�3�Θ�g��s�����ܹs���3�jE�n��2/��͉B���,/�\�r��7oppp��p���6;�#Fۻlo�(�����C�%!xZ�6�����\�y��׮��=d���jw�����mc3K]V�'�rAUV���[���-z]��=�=`���pk��ΈN�+X��(m�V�n���p���=���~���6���p���>���ӓ.]Q�JZ�6[[[\���kW��ۣ������u{�[l��ԡf�*9;9&��d�A��	eZ�Y)*������p||B*ZM�==����B|s"����#L]���ϵkW�rp�������sAPZ
�ҫ�r�d�������z<y��?�=z�d:�p�+��7��Z�7��x��uD�}��Y�HV�{a�Ġ�� �	i������ �؈��b��k�����B|=V�F"Q��b�/��Fr���٪��o�zr���� ��h16`�!��)4A{�/[kQ�\�[ ��$�քNĈwNZ��㉍��^8��_�=ew�����o�������cB@�O#:J���QQ�� �6�x�$��(��Q���8��B�+���*��>�����~�!O���l�SOd�I�)=�C����Ʃ��(�\�������2�N�^������*�hu:��\B�)lk���j�>=��?���=E�C��|����I���6Z��BEaڴ������7��D#�@k9�`9]r:>���ǔ��<�΀�����6�v�Vf%T�?FG��P�%����'O�L,Wc���v�~�:���	��rW��3�O8?���#�r������mgow��5�������g6srz�l��*�ʊ��{{�\98��iK\��~��آ(�����x�����Ea0�2_Γ��2��fw[ "�����Cl&y��"������/$16�zT�U�]`�������ի����E!9W/�UU2���SD6B�4�7"�bca�cM0gMk2�G��<y��dBH��_Fq��ڭ��ŪmbN/����ȴ�|���o�iZH�E+�	�?�F1A��'��5A*�%zq�Ù�ɰC�^ᵥɯ>W�yY�g}�[I��Xb*-n��JA�hR�W4Ѣ��{1��`/^CsJ��c"!(� ����j���*A�)����N���~�F|���+;�����(���eV�H!�ȇc�����~���yF�HA�GX�-������d���������Ɲ;w8zz��2�1�fs�x>��֨���,���5�Z/�(��2���еEr�l�R���u�t�]Q����*WԵ��+V�
�4&�k��ל1_Ftj���:Դ��:M�k�n��2�`O&�hc�'<����&�(���=݁�b0���(֩���9��ɘ�rE�VX�f8���M��$�F"`N�9��l���)}���elu���=����h#��$%:�LX.,�
_UTN�F�!����ۂљ�BK�����r�`<�1�N��������L�S�jEUGZ-C���t���-�����\����G��п��_JDq*Y.$�TU�)ZtZ��=	��e�l6����
����"M��M�	��9Ĕ_s��tFY��U��k��(z�Zq��<{Ϻ/��vG���>�u��Yh�O�h"�íHξ��T_J.����&��������|N
:�����~\�f�ҵ�%��7��O���M��7x��o�B�URZ)��A�Q�*BB��*�����R|�:�8SZ!�:'d���>)����裏8>>�P��*�I��\:��DʉQJ�q�6'+2B���t�����\��&޸�O�ף��^*��} 7�V�E��D���W��uD#�c]�ؖEGijt��1����h�
8'�����\�aj;�.�@�y�(	��
����I{Y/H:���{�����HN�h�|6��v�!&����)�L��lC�
²Z⽇�Y&�����^T�K��d����EhB�ӡ�j	i*�_,� �I�'dnB"���yq����ĳ����/P��"S��W�	>��;|P�J~v>���CV�uhW\�!Ky������#>��Mbf�Qd�oT���_�8������Ϗ�|S����⦗A�@��ۼl��F���������k���<��+�!&6������>|̕+���~�o��_���ާ�*(�RJ���A{�r�C)�J��p�ҔSUD��ػ(4%
�	�)�w5DM�nQ;�O>�	��?5��8qLJ����r�)�ǖ���t;���q��4�s%��J.n��@,���O�ק��-H)��B�^�dC�Xu��z�����B�a2>��@P�L��L*���א���T�U�b1_��`�F-�Y���1J돋����*�Wy�`E�照0W�~|dQU�+�T���*�Z�u-���0:#&��"ϩ]MYz	�h����rI�բ��Jq���5F`�^��9o%=a>���D�w��$��RU���ی��Y�%��,���׼`c��a�/��R��QZBpu]����$�e)a�ӳ3��$��n��đ���\����Z��E"V$��!��_}�_+ί嗑/�8��4�3EA�y->|��+W�\R�E�S�%*B�)���&�ǈ��� �)*�mNS�إ�$)���TZ`ҴҸr��j����O׊�c�����F��3��h���]�]���F J3�k�[i�D,�N�C�ݦ��C�!
��l<���a§U(YU�)��y��l(N�3N�[����!EQ��2($���U����rFYV�d���F�y�E�e�>Un���Y-�,��*�.(
����V�h4��w���.1*H����1	�KQ�|�ґ<+h�9y�Ū,�OƔ��=k����pg��h�x6�\�,���(Z��.[�>6�%ĈQ�� ����cf���c4����V�Ea��W�ı��u�\2�Ny��)!�1�3S�T�7��slmm���E�ݡ��(+�j�U�j�d����fUB��ͦ4�3��h�6��jŽ�����x6J �Zq~-6�+�8����z�q~��UP-h16��Jx3����})���NU�uL�U�I%\+j�+���H�jS;ǟ�C�oNqJq��/|�[������o���(�ZS�:U~�񢛣@���g�'�y.N��c���?�_��rrrF]�0Y.�_����E�Y���x��h�Q[�5���4�r,�K�N�999����Lg��^����.�~�V�M�8�/�ܿ��ل�b�����g��:��n��׮R�jNNO8=;�,K����������)˒���>f1Y0�������)OON8=:�+�TF����w�7�sxx���9��s���ls��U�]���3��,��yf���K���<=:����Nw���!{{�Q�E�V� &�)�K�����O*�o��KՁf��qsq�	Q(���(lcr�^=୷��{����Yf���pw���ij�׹�º�ps�7�'1JM���1���c�|�1�=�^ܨ$4����_+ί嗑_Q��Mڭ�ŪD�Ha��ic���)�M��.��to��\
�
�q�(��5E�M]��ɥ��S�J��������?���#>0��T�3�ƢH��i��HS��1
Xx���'?�w�w���]ΧSrk�|�/Y��Z��8��P�CMn���{lmm���|r�s�آ1�<��i㪊��c=|D]�chu
:�>�v�V�bggG�c}��?�9�g�L�S��dZ����N������6�jɓ�O8<:���:�ﴹr�*��.������}JW��tܺuk-�ق{�>c�Xb����U�vv����]�ON8�NQ�3��fw��pH��,EY"�y����t�|���=}���SZ����t��,K|�YZ k� 0�����'?g2�\,֊U7 �I��=��jO�ƒ��sn����ַ������^�Z��D16�صJ��?j� n�9�LWN�������ƿ��ɧ?���It������Z~y^��Ay����?�N��z\�v�[7o�=���u���(l�x����_-��� ��׽�#@ɩ<gmق ���˅���1w?������}iOmc��|V��w����.?���n�=��א���ᐭ�����`8d��Űߧ����'p0�����z�z=���� k��{pzv�r�DE�K��˜��J�Y��Z�`l�e4����*�2�L�ϗ,sB�Ȳ�^��j�b2�P�ej�����Kʺ��~rr�|��\,��FK�,upYN��bwoW�Lfs�˙T������ွ�=��̦SNNO��1��m��.�n��|.0wJs��u���9>9a1�S�%.a�*XW�N�S橧q�X�|I��t�}��g,ʒ�l&J��c9��X�X���fҗ�Z.���f9�^��|FU׬B���%-�/7O_-R��(B��Y�����۷o���mvwv����t;O��/��G�skk�`0�����_�+�?90~-�9��_}�����ޡ�����k��Ҹ?�(��-M���p�"���k�q>wi������+�"V���ҫ4X��L�6��Y����4�%��2#�q�6��,e�b�\�\��+ʪ�jF]SWu"��W�Tu�O-������.�PY��U�V!��:�J�DozC�"q�	wR��9f���ç<x����r~2c�X�g:�0��=բ��J��)ggg���3�LX�+2#��4}bV��T��K�J]Ղ@�XQ-�8������+��+qc�>1V+i�_�V�#F���یvF����?����Rz@3��V+N��y��1�=�����c�����G��c|Y�v�w-K��]L����?y£'Ox��1�>��?����c����:~��xno�~F"�k��b�&��1��*+���jI�Z��tU�~�Q�2�^Ϫ�pU�� �/ˌE٦��k�Z�ZQ)�����V��eř~�d4��E�ߣ���?HȜ�Qk�E�Cak���N��ԩA���Z�+�j_-p�ϙh��]Z���b�4��i��9X�E��+�!�̹�}�{�Հ<+)� ��R�3M����
���fgk,ʂFQyOt&3d�<�0�`�%�#B9%�TЉ%j �N���-�rL���=dow��k��=L& ւ%�Q*���z��x��眝3��p�w@�Zqvv���)�r��Q��Z�a�Q�%�"���F;t{=�1�����ʈFxS;yNѓ>ҭY��RXe1:�������,!46�s,�D�<��� z��6��K@_����l�:��z>x��I�����Ȧ�|�Ѽ��b�^V�i$�#�5!*��,XC�!FK0����2Dm�FHDe��ϴD#�AQ����l@�Q����q����b*����*�j2��]I8D��_���d=�ϋ�WJID��(�q�h�U$�oB$�)Z�$����i�r�8G3T����tQ�ߚ٢c��p�uKCTm51�cR�.
��Ӡ����:l���[\��R���	�!���t���y.��;�,�K&�9��3��e�<Q&%�ΨQQ����^��`ؿhc�*i�W
cDф���t���fggG�Ȯ���he9.a�z���R;�F��RJ
�"�r�M3D�N��Z�/0�ժ��L��S�8�"�?+�k�Z�4��u��.��)/��l�O��=�G�ѧ���1k2��� U�Z���D-3F[��~Ic�X��jFTVZ�(y��T�A4�8����Z�H��\�⤗�RH����Tʯ$���n|w�<d�4�f��^M(+����$5���on�X��KP8_����X��-r#��Ps�(�*�m�Q���h	�6�-�I��+���ņ�A6v�ĳ��E�O��F+PA����r�cĶ3L�5��d<s||JU�dYF��a6���/���(
:�L)�|��-�ֆ���V�f4�����v��b�t2a1���&�9�9���kW��_��|�;��/�������}��o������N�̈́B����fEAD�\.p��(a�Q�@͘J��������*)c6��Ƹ���p�J^�e5kW��~~?�_���ǟ���%�j���>{*�f�Z��4׳4�Q���2��%eUa���U`�%�s�!$��к�f��O��Z�}n�y>[[�6)/�J^LDkA��z�҉0�#(Z
�����P4!] )�����T]��uEUy\��O�?�����X�� Ƅ1���T��ob��f������r�T����{���m��\g������ٜR�_��Q'"X�PC�kJ
�eZ�t�t:a&�r��֓=^<n�e�JE��<��cp���4/�R_|��b��[BD�rH���(�ww�r�
ׯߔ
އyp�!���:t�XxQ<Z;f���'O���̦S&��傺�����^'����6��C�>��Є�A&|�Q}2�݈.oJ��Fs�'jt�%���Y�@�5��r�aM����iž��#zO�n-~�HNP�=1xa�jh�|�+��H��A0=��1�y��}�������|�1}�!w���·w�����Ï���>��|�!~x�?��?� �|~|�~�~�!?��|��|���䃟��?�)�3��qu-��X�:����	_�!��w)wt*�WBT+a�~Z�.�z#����S�MHc�P�4�Һ	�6Δ��n˛��<#��4[�;;;���1�ݦ�)�/�����O�Ǔ��E���!�UA�F�mu���tr�Z+}�ؤIĻ*h���������E)��̄�h��ZB��R	�Od��1dy.�P�$��7)�!+
F[[��1�8??������c�����P�t1#.hf�	O��9z����c�>}��|L]�Bnl�4��{!Q2}%�.9�T�/��+%U�k�g^������u.3J8z���5�^$͚}V��^���b��l���_��5���|����0��y)�r�Xm�~���~<;;'39;{;�z��c�Z�4��1J�������{���T�J>Ч�cģY-W���1��Y�j��J~�%���D�b܍�Ai~�?�?�������Y#�Đ�JC�?�7�{a���|�`�����i���*��������������ɋ�����H�@��4�h�U�UUc3M+/�}���>:h>�.kb�t�}\Y2��XΧ,ˊzY�����W:�PS��XGn�s���F�-��_���ΐN����O�<����4�V�����\-�������t{z�.�����h�{�M������g�����,WKڝ.���C�V��'��<}�EY�iM�eTu-��9t�Ӳ�����[o	��1��O�b:fU�k6y�e��Ӻ��1Pm������?r�����}>��c&�g�K��h�D�{����$��W��j��g�/�������}��_�kloo�e��F� �����5��wB:���D���ӵ�w����C~��]>��#l�ZC^���@����Sgbk��3M�&+0Vb3�,�u����I���8B�"n�q��j�Bo�q�DYV�n��u�~]�TuM���t�d<a|~��x��(τ�����������x�d2f2�0��O��'�4�/��|�X~?������|�sAr�Q�XX+�g.�+��Z�������;|�{ߓP���]�TU���5j3���	���� �0W�����Zq��#>����NXT%E�@^p쿈��0�m��X�TS�ڰ��Oar�Ւ��G,3�z�b��2�L��2�[�*�w��R��v�w�u���ɔ�;��-:̗&�\�0:'�-;���l|FQ�h�m�<��ш�̇�sT8G�bk�g������Ō�d�d>g���{OY��	�h�d#r���EA+����FY�b>����W1y����*�%!jJAYה��vK
�NOϨ��D��!`�p~�`&7�_�����f��ׯcS�r媢�W���k��.�!d^׮&��`�=u����	��k\�89=��?��?����x�� I|��Ӥ>NQ� ��Fi��>N����>ί�+��#P�~��3���MR� ���9����}�g���b�|1g�h����gSsi(_�B|�\.Y-�̖KV��e�/Y.W�W%e) �Պeb�/W�x����S)i�|�x��	1������׮]c>�3�99>���lm(���OO�k�`2�0�LO��g�����b�b�`<�p��=>��3N�N���V�����~��R�d�h J ��Q*�d�����,�KNO��N�u�����l!Q�b�%x/�"�H�Kn��٥�m��9�O�����`H�n���9���@fyQ0�|`�X�jw�
C����mwn��3�L��f�U�҆�����ew��`4���'B�<�31	wv�X��Kye����%$o��F�����',�
���ak������`f��&j�V
k4�x���ONYV+1�PĔ��&e�f�,VQTދih�Yp�C��,�&�)��g����Nd�ی�D�%��2�ŀ=g:���;�q��}��~�G�1�-ċҦ"-*��ˊ�Cf���lDi�V�k������+gJ]2U*��2���v�/Wx�iwZ������)��7rQ4�X�i
�Z��%�����F�l��
��dބ��X��4��[7o�o|����E@UV��ɫ�����Xw��!�s	�&�;c��<y$���c*_�����^�a_R��n�jAG%��MNE����w�K����䔻w�2��R�"F��e����dY��j0қy��u�#ڽ.�>�K^X��m�R=9�{w��k3���۴���b��9�*��<y�v�����9=9���'<����jI��3�x睷�F8Ws����)�9���7��PZ�ӟ~�trN�*l�	�P��Zz��n��h�j��|HUU�Z
�q(��@iic���4[�h�Z�	���v���a4��'�0>?g2]����'EQ\T��IQ	r�M��ʨ�߿�իܾ}�VK�V��G�<�f�6�Ԭ���J��"��==�G?��?b<���x�J@=^G6C�[[#�EA�g4k�
�^�Ƚ�C�_˟��2T����7B�AkY��{=���N\.%d�j��J����$��i1�%�
�g��QJ��&\c��$)fu�
������6��6��{)w�k������|f]*�?آ�8�Bk�
�%��3��%�l�l _^�W�9N��tf��w������<x���|	
1Zy�V�����\��
z�.��6�^�v���v�M�����LY���Ʉ'GOx��!����N���~�����FcS��|L�紊6����C��+O��a{��o��֊�d��{�X��D"W��we�����gg�,�31^��]�5y�C��筛�ɲ.�rʇ?���Zb���x�@a3�����^��̈́��U�p��k���v��>�s��b�[�(]�Z���ԩ��M�J��E��Ġ�[�ڂn��hk$������kV���`�_�������o��ش!��u]�X.9|��r�,o*�Z��J.)��$��Zq~-�z��2V�f�����v��r��*+���C(� �c� ��/}�(M�(�W{�r��4�;�1bn(i7�(�_V.,o�4���\���𤘆M<�F$����M8�]�B��*�t���Fg���_�D�Hq�%��������1p>s�䈺.���+����WLԠ,�Ռ"����~��ርA��|Q��W��0��srr�����"��s��Mvvv�m	�A2j��$������09?���tl��~�U�89>���S�#3�~�go���==:�l|�t:�*%�Z�p�<���w�z���Tˊ��	uU�#�CAG�hg���=��C�\� +�EYU�ڱ��>��j��uU�b*,��7^�R�6ji2��Wb�PcL!PG��0�<}z�jYh� \Ę�*2�TL��i�G�N�� �Ͱ�J?D�x�^����s*�ׯ���y�w�UU�cH},!(�z��������%n�Z!�(VqHʊH�����7�8	!lĶ��Fk� u4�jz:S��d��F�G���1�%j�%�XI1J�5���X_�85&J��
R,����AQ����	*8bPtRR�
�(�|>��sZ�.�NO�ѹ ��ͤ%��jUQ-��WV�%�{TT��t:��6Fb�ԾN�R�}r~�j�b�\�eV"!���Ҥ-Y-g�h�k������޳Z
X��s@�[�R�v��`4�)��ӣc�J��!F��nަ3��.
!k��B����
��9���;)�q!b,�v{З��Ћ����r�SǊXk\t+�,�K��9O�R�+|0��F� DQ�Zr�M
q����ncL�DV�i%!�Nyr�`�|�8�m����efm�ZI���_�7�8����bN�����FД�%�	�x��ڗI�8�&�7��`M��(9�7�UR	B3e��*+�12�����C��Y�a�i��4�{��F#�F�hd�JO�S������3�SoBd�N�3�⌀A���zr�Be5�圐(�6jA
&b��B+��!79�< �Ar�$�'�1B-L%F��9��d6C[����6dZ��Jj�*�AE)S$�'�U-=�֢C �b�JyXU��SB�&�̢4-[��U��DPFº0IYD�Q$������oR̻�GH$y 8/БM/�7�_N���(�*�YT�}�`G�px����x���C��
�#Yf֍��J֔�l�Yc���u�P�,����/#_^q��ɫg|�����-I�fW�_���l^K�t��>��}���ŗ}���e��y�9�qT�:񞪮Eq^9����UI��D���t�m��������o�h�>?��l�Y+NY�F%��T�KI�!QYf3��㱺���%H7Hc쳋7����.[�[}	���j�#Tiױ٦e���f�e$mbk9�\)�{s1�� �[#0{e�����h+�a�	�	��
)�QJ±�]x�R�)�9D�s��dh+f���B���K��P�� 8�J��V�䑢�*t�P���/ش\��
$3�ie1�Fk�E��ֶ�]%HDQ��31�S��JaX�c/�sH��N��M�:���_�:~рS
��V�%�S�s��k-=��E��	O�<aU�D/��B��z�R0& �f}��HƳ��K�0z_%�8;Iqn�Zq�Z�
�����%Q�4M�����K��vIJ�h������|�4�3lx�IyF����^D������׿L��s^Wt0h��kV3i;S@S����^����~]�xW��>��5y��#m��Y�L��GQ�z�q!Ĉ2�&���WI\W�F|TD�sE] !W��֤�1�Z�����RQ�)E�=uUA�(-yG!RL����	[&�;%ׇ�0w�\���V	%9F��Oe��Q�ѣ��PWK��E�\M�����ߒW���f5W$�L$VHb�V�����Jӭ�Qw����8�3�����~��G���Z�fW��Z��,���	 ��m������Z�G��2_&ߗ���annnv��kwq�5v��
_�� ����N�,��%N({%�^_8\���v���SH���ۡSv�]ph%Ω6��-�����ḩq1�������1%�����nW���D��u�fF)JGBL�4���fu��DEA�	�Żu�(E���tB4Q
UUj�H�I3R" N%��,�yٜ��ss�
�7;�����&1Ј��:�b��C����)��l�IU���C�5�jr��M��L������F@稈��"1o�(��Rr��	z�{���ei�"��I�v �$�)���a�ݠ�;�5���5-��H���C���u���9i�ӭe���;iI��$~O*�"��=�Џ^��H�И]��������p�z������ԓ-*=�=ӛF�iBMQx�sH���n���L��GJ$b���V�p䎼��%Z6ϩ��I��J$�ኅp˫��,q�!ι٪9&��䛵� $�Ƅ'��������S�L,�x ��JU����Գ�,"�uC]W4M���R�h�Jz1i��7��IN-=�J��h�]	V�(]IQt�ST�E�Pf����Q]4RT�%�t��E]	�1��5�IM���PxM�5�Q��bޢOײ��I	'*��p�ᜧ#���{b]SǨ�#��\G��{��!4T�"�5e���v�t:&9����!Z��6�����pF0̵���]��$� Q3���gD 1%>���-�����fU�A#�z�cL��܀�(�]�eiFe�<4�>W��8&��H#D��l<���͵kW5��-��Ł�����*CDeVF0Er�J���p$�v��}�l�SHak�Dv�Z�}�>�RV"!xDۃ�:�lF>�=;i |����R]��4���:6�*Z�Z"H�y�ڧ["�ǌp��<#�"'[��Ho\�-�3��LJ���C�?��ӆ���-���{��7���T�H�nt�7Mc6� gAW��)g;�v��L�#Ĭ[�eD"!�!+�����^>y��fÄ�I�"�H��8[�c�#3N����lln���J�<�((R���yh:�>.%������!uc�(lŝSw�ŵ���r�pN&�{{t��5��g4����Dkp�)NH��9'��c$�
I���U���.��T�C�6���1�h@�����E�Rh1��!��:��XIʤ�X�T�:L�H��eG�Qp�X�+o'����qBl��{�+
����?����~E�f�4Ī҅����]z�)F��Q��bQ�%�ނ�#�st�&C ��|_Ӕl��Y=�HbTU�"'x4'�t>�B0/�|�P�po���6׮]���Vu'3��0n{�b� �t��}��|�Qp/ƙL��M��(
J�>��1\Xp*����m����$�4�� �W;�=���� �����־][ �H*�BZǒo�Q���*���l�q��;M�<w<G���|]6�r�}�^�A�<��1>/j�ޫ��
$0�\'����x�y����e����9�(ͩ1e�aH�`�p��E"��ńÌ"��D��ɓlnn�������I����ʲ{MH$]e@T��i��.�\�F����;�[�����XXJZ��X`A�����}?�w�=����<��9�u���L�}1X�ZW�i��c"O>��g9�ۅIG_��o�5hsf(˶�~�
�4�4o̹��ʢ��?#��Z��w�=��z5�Q*���Ρ��hI���6ER<B�3$�8�����"�W,}B��^�'���m��ݣ�x�.�a%�w@yt�����Ԧ�V�yq�E��Í|�}���^��;�/+B�U��L������:U�,-C���Ԏ*�d��/"�=�	�HI����*q]��V����������§7��w;NM�+w�%�kC��K-�}cW o�j�߯�,���h[��UB�BKP��"�oЕ��� >�� Xڃ�'_�h�}��|�to0���]N�~��ZO�ɶ���{_H�� ;}BLۘ"��8����X�'#��Γ�Er+!U	���ؿ�����u��ƛ E�]d4� Aq�ѓZ�N����$� �v�$5�L�Ҋb,c��L�	�E���݄�7g��+ǉO>�z��p)�3L?o����L-;���W[�y\c���2�5O"�f_SE��J5_���C��]��j�W�w��Q?9����ɝm�ْ��)lZ���⟾�E�L���*���stt��!�!����X�=�׋�׷�\~�t8$a�Y��~< zX#�wB���̰��K��ۍ�p��! ĳ�<��#��C�}3���[:���>r���6�ެ�ݍ0�0�(�>���C3�=q��vN�mƽ6�����	�:������J��t�0s�^����G�<6EUY9H-ߩg�P�/mʊ�19v���w<���~��B3|\b����I%#UO�8�Uf��8���at6��ȓ���s%�峊�qsW~q�2a��\-�ߩUo�"�v���'�q�p�����c����^
	�vWj�SR+ww����&��ZJ�?��#G�CL\���ʃ�?����ҥJ>>��:�S����9� Z?���~����/�t�=9\�t��1�=U�B�'��Pq��y��;����};_���{�u��K���w��;k���Q��+/��B�9u�;Z�!ޜ�4��:����Q����QKp���LX՛GN<������;?�;��24{U��8�@�r���ӖS���=��&���3��կԯA�z9uu�������`L��5^J�f���%̗J�Ŀ�<Hڸ
c�]<_{>F}���L��
Yߓ��9���+c����{�}��l�{Lc�q?C, �:`�c��ٶ���� �]���C��i��y��F�����Y��Ʌ����v��8��ü��螿�CK�([��R�O
���oǧ�έ����j������ʓ����/�/�9��A��	@%5�������MW��@���jP!:t�<v|�@�����F�&���ۏ�~8��c:�)z�x��qN�qI��~Z#zɝ�K������mS�§��<�����=B[NF?�.v>�.?<y��O"�W�t��c�.b�����'�<�Q;��ϝ�w,�w��Ϋ�Q?��Ӻ�����T��DQ�,l��46���u�~}sp��4�|�܍h]Ӎ^Nq&���cѩ*!m5/}r�gɓÂ[�Ե�����~��S'қ=\�>�����s��n6��o�f�����=!.}R�Ǎ'���	ʦ����ZZ�G�<���sV)�X��#�b���B_�H{6ݤ4C+X���7�f������\�8��'M[��gZ5��M�X9�B-f�s��'��U����3�<#��in9\ʸ�n<�ZIU��)�8�����S�o�C�%�/"�B��P-Y�LR	�Z��C��lW���a�9�����8�d��fVC��~����P^��aUR�/>����VN��q9C����s	Ml����	�a���8v����]{$��������']^�����7yEFEaj���c�T_�^Z$� ��%�`m�)���������I���8d����F�ڥ\����B�Jv���X��FΟk��P�>q�Fr�C\��㮀(���K��syARy���`K�&�w�s}Ghm�4���������g�����ju��ǌ�^N8�Z9um�G^���z��E�������]��G�N�z?��������(\s�<�p��ߘn��9ɇ��.�o���	F���c�Jpm��U6e~�*[�+c��� �!���#Gf1�E*�{�%E�ռ�J롌�3fw^�\Y�����TAh�T��^p�j-�F
Uj��/�BˣDf��OVP,c ����0ʸ�%4ya�
6�!�6��||���������m��l�je��΢�	@R��nN<*��\A��p,c[`w�j삖2�~�g����C����B(�͕��j��8���u��D��@������km���nn��i��Z�ޗ'�L5[���E�M���k�.����F��}���Ӏ�Y*�T\Ir �%>)����'d�ϫ�鍩=���N���i�G�H�r����z��.<]ےf~�����m���8�_;��ʠ�_��b�Vr�v�ER_�\дM�K���L��¤�tEf�pIE��)B��l��6�ߖ{�l��-�L�Q֢�D�T �ql��7�'�v0�/��Σ���i?��\bKd�4���V�#�%7rK�`���ܻ���4P�$1p�B�h��DE8��h��_�L�d�[���2�2P��Y�Σ�[���@��a��L��:'��[��%,Kg��K���k<�E�YQ-���;�_�R�%Ά��:8m��ݜ���O]��h>O�e_5�I���Yꐥ0�-���~9��2X�F����w�IbF��Na�	]�Z_���U!�j���DN.H���:���Mt���q�)s�4�	��ۚ5Â���4:L�Z� X覓�9ө���-Hy�9&�_Q�5���m��C�ҩ�dH�}�}��3\�n��	u�T7_�.~CR"݆���JBN~=.0�	�>5�M�$Z�ĕ��'J|~��G}L~�C���Q�{H�*0���y.����k˷�Tzz�vn.�8����Qd�B���Y�������{5��xR
�E6�b��>�.��=��;{���z�0FgI)S����$i.�Goⷪ
`]:zLvܨoͥ�u �Ҥ�c���6K��1�N�����	�g�g~����ڀH��T%櫐�Z�r��M*����v.�����S�rt.����ۑ�-�@&�1wܠB"����s�s���y��s����H�:W�>���\���k��/LaZs�ZF5*)�ϵ>�\����?��_��3��|Ʌ��w��o�ͳ ��<9���;�â�O�Iu+�+$jW��"�woPXDP���>�,��<�!Bf�=K�_@�u'ID��f���O0���?۰Z�z�V�Mu�b����������Ws�v�!GA�"�(�~�Y�a(@;$~���./c� ��W�[[[#e$�N�α��{?�#�C_Lz�	j��E�<A~E��e�2)�;U����,'��>^�V^��Nӹ��r-!2�ȕ�[[��C�1��li\��eI͂��=u��nUR
�ͨ@>��FF:�P8�w]^r�\=�'0��۶�}̇����v�����_�t��>�H�9���a��/��4�.��w�����V��m�؃�����%L�5d��a,�^�`���1���f̣�g%����s5��v���[��S��nB1 ����@Zv�"V[��gǕ5����3��>Հ3M��k�qQ�,G����g�'�v��}���f>_gB/!+���+[��c����7��O���w��/��U1J'��.�y������l&[�y��	�SO����[��m�ؓ��y��C� Zr��VQ�;�?�(ه��������s�����h�3P���W}m��b�|}9y��_�L{vö���'���@ʓ+��A��[��3ˀ�����Iʋ��e挳eoq���=�/��!��7�O���/\lzeg�{��1������c���1�v�y��Ǫ(h*�'G�s�9��`��v^�E{�#��w�)?�P�k��l�����Ja�k	���۽��@n0P�����t��ۭv��+���?��5@#�_I`D����T���ܚ�����:N��0%,� ��������=��w�_'ٮ����e0�'&.��D�Px[na�\�D��&�L&,2
�k����~�Q�'?����}V�`o� ���+����U��:T��m��7ٍ�����˕ǠT���x�q[�/Z������ �	�f�X%����������+/��y�眢rX�wz�+��ܥxOMSQU��Z�����T!��E� ]���
�������,,Ǆ�ʈ���r��ae����-'G��W	�ܥ�CS�P��mq�*�4����%>����uio"U�������f�G�����1S˱�����:���й,�A}ķ�G����ZB����GH��1�+���f�Ύ��M,|��5C���gq�����ҁȱ��ݤ�^Y^G�c�"�i<�E�t��l�+�Ѹx�u��������*��u�n�E�1b(-�9�$K���b��E�h���m��F9U�>�:�����u��9�t�����	;ݞ���~��DY~��F7�D��O[��}N�����viĞ&cД��LZ��|��e(lj�ʰ�ʸ^���9�
�
E�z/��)�����W꼰��'�����-KE�^�ِBv�xvR��m9�Ŝw��=�6j���Ry9��b�B,�j��.|�F�,,,�,vv�MP��9Sǆ��Y�9G��#�;����f <~�=�e����t�Ƌ�k��ʊ��&��K{󤮅�,/�+��������H��#�^�\����O��le�R�����`�R?~�M��q��� ��ky �����������CysX�Dp���b��.	�$w������.�A���c��;�^����s�M���N�q��_%g���i�d��2kk�ߎb����W�4��$���b�?��݂�jGe�ʧ�fc�����������T%�HY�Q��I��e��U�5��U��W.�+��N��}�&�$��b���������G���p�D������&>>镕 w�<|ᛥmh{&�!��.��ISN3@�Vy���t!M�ށ�(�K�CԚq�ʦiL	�S�x�b�������GC]���U�e����c��v����s�r��@ð�",�Xμ*�=	�_Y^�x�}��2w(��R`�D�{���u� g��:���ϥ��ӗ�.S���f)s�Ch�d*-ܬ&�'��W��H�nX�+LA(��[���mQ��-�w�WH�UX�O��˰���=lC/s q�/,�xx��7A��急B0���T:��Љ���쨶�����'TD-u��^�_n�PQu�7�߯��ؿ�i�߷��k仆v/,�ئ�x���v�p���t�
ǊzhU٤�|����������N�.��3����aQ7U�9�۹`j�ilo�9�˧�SYQ[[;e��>,�b׮��Z�������챍M[	�g�{�p�LY��k%\���N�c{���n��sI�U/@f_7���Ԟ���´��3���3�����Z��?}\7�_��g��յ�l�;�����rO<>�^�X�Ziw�*�^3}�
�DL����� lL❝�y�> C{�R��'2���uB��U�	�p���)��}��'~����7}H٣~o��]���"�
�6_}?�
E�
tya���*ՠ�=�E��ywȜ��ۧH����n85����&�pޝ�7h�N���{&�n�ѻ9�C��!O��]�5����m�c����|9D��t������ZO�r�?���7nB�nO���d5�P�p�,|��f�L��Y�"��6�����	5e;G{��~�*����E�yB��Um�8�
̟�y98�
(�RIs�#����7����E����?;'�-Ɉ&&��j��fO�0��K^B,�p�Ʃ�7Jl��8�,f6-���C����_f���"Z펏�I��e�3�z7z�ާZ��/..�y%��9Դ���&��y�e�tH�<3�ɧ�������J@6��.��pEv��3�F�wS1�m	���>������2T��m��Yr�oM��f�{�/�0���t("kKBYMǦB?6TTU�"�m��
�ҳ���a����{��Kzv�=*WA�cE)@����X_o���6�p�}�Xs��}�,o�H�g�<�e�˭�_v^�p��)�7o�
3�OH��d�iȋZ��'�DyZ|��gl%o4>��:?����
�`C�5��*F8|�X�y�D��K���WD]H�G�~�WY�\D���j�$V9_����1��VФ1s'l����5۫��[p�dZ�k`�E�m�?j�����*�7��JC}�zI�OB�@�E�}��f�畁��O�Z��0ƣ�f��J(9���ya�ĕ�k�!}�j:4��@L����S?1�CN��l)+�p�L �WP c,	 ���L�Hq�J���V#V\��̙;ƄN��P�qFRx�,�cg�F� fܤ�:|H�C��	�_�g,Kk��i�fԔ�# �	#��=�������Q�ʢˡ&�<�Z{3��Y���Wr6A	�C�I�sn�x�}aʄ٩��q%��	ܻEU/J�����$����6���._�nD+/%�_�4�����1����y� ��3'MI����:�T�������2����rr����zڊ��4�#Z��`���y2jaw��	Vt�߰X�������6P��c7 �m����A��h��ۣ��\h<'ig=M�������26��0�-v\L#�l<�i��F݄2%�'t��sN�����3�T���3��6�8y!����q
Gh�i�[��s��NU�_�7#L��+�n������n�`%�U[2�+'L��N�b无��[Ir2��o�����qH	�4R].J:����{� I��v�<~C�8V��dE�NJ�6/��1�?����}�k�{E��	F����}��ꄢY�jo	��VZ�6Z­�	��0D�ڐ����S
'&EL�����L���J����3��h�L�":J���3I2$�P�����)�N��w��|eXɀl�OJM43��%������}47�����/h��V�#~&LV�1��n@k�ENE�"���#�7���KU������y�p舺�B�µ�,N�mаrѢ�TU#iՠ��}�Œ~~���ۢw�K^%��IF����^����.�)�6!�%�`H�����U�;nAӿ}�,�.Ơ��nH��,�3�4L�yJ��]����`
���-�W���������G��e�r(����'3F=Z0x�vj"��+@|�� M��������	MޔNN�ᝡ U�W��̾�#� RT�.2]�m����2O,,mtK�ɜ�����Y����hSNڵM~d}t�LO�&Õ��/2���#��5����d�[+T����N>_�Z���R�P2�If�=��72~���n;��h��_�@�c�b����$6O�sE蒧{՛bY�rʃ�W~Pb�9���ɧ"��ᰰ�+��G"�`y��3?:ޱ�۶T*=�łݪ���mm���
x6	��D��E*��D�����5�+R���n�������$�>����GS�!��C��g�4Df2���^Vɚ�k��j��|q�z
g
�_+g�^��C�[�l�,B�;#�M��g�o�����9��f"<�}+ֈ(��<�x�	��nL���$J�f�7&��h>���NnB6��y�9�"�֐,/f��e���\��c�L�jPNr��4c�W��I
^���R܎���kz�7}�4�L�Fu��ҧ�^O"�l=~ʨg�=��_�q��-�")ɾ2F#��r��u7U����9h���os�E�Q�E�9��7z�y{���UE�g�t�XQ,5B���v�*I5�6����20K:E�.�md��������^��/!����D;.o�c��G}y��x�L_����D�ʥ�k�'�(��C#�e2z*<sjH�ŭ�ۑ�C�m��*��̟���՚���H�y�zmlO�n����։N4�6!Oz��?�${�o� �~k򁓄���E���|d�a�&��5.��}c��P��^�O�!�O�rݲi�1�9��f�c�ӧ�+�7�U�Uʚ�ble��6���t��'���-�E��*��b�)&C%W��w"���J���Q����[q��:�o��Sm�L2���	�l�㝬��8Ns��T��"I5��|����fu��I���mp��ѐ��審���H�Obs�/FR>eeWn���3�������_��n'-�%)����IX����]'�5���qb*턻:��o~y��M`>v���K?�v'8(�Cvj�����g�������Ig�V��|U��jJ��O���.Q�h�����>�zu�R��)1�4��TCE:1[��G�g&:SZ��R�B��%`�8d��R��1%x����5;���.�׍�*�	�Qu^��ϊ�R�iyӣׂ��	�Q-�F&T�m����I��s��)�G廦�U�A���#��>L3�Ҋ��2yrShݍġ�0`��ֿ)����S�p�$R��ƛ� ����3����c�� /�d��
$:��B
a�����F+M����g��m "]Z\_'���_(���<�b�W4|n,�3����D�CqX/|j�gI�A	-	p�;,�]�Y��v���D�7`�ޞ�F#�����z"���m-=W,����+$&m�2���"p�N�#8 ���t�gT�0,��s�s�כ��F|����F}y2�$�#�.��O;�a1-\'�S��Br�z`Y�����w[V�+�8ܒ��lR�f�ь��G�@B���+u�/l�.��w˄<|DDէ56�Hc��V�r����N�c/_J^���{�@8RW���s��>~v1���Fl5Tcat��#�6�&$ڒN:i�O� !_4"��8�Q����-9O=Q^&�Q.���̫ޯ�v]�&�0ű���m�o:�Pwy��PF���}_|Q�"�`�^�]��z��/�W�^hq�,$�X,(l7U.�*��U���D�Eve+0�6-����jM�����_����Z��'蕋�ɱ	�S���l��5*p�K���li{K6�d ���&j���S�u��y~e~�����b���HP�
�^
x�T௨�m�����
	��"\��3�]���O�}��u�j�R
�� O�T�eU}�rfI4Lx!�ٱ�z�wø@�#1��.<$����n�k,[l|[�Y��a��|���4�H��r�
�(f$d�DhzN͉�D�+Q�&&b]da�Q��ٽ*�\3����f�j�P��z�(��kY��|Ce���!��atw���gE	�M�-#�k�ga�q�5�ݷ�GO�ء�J^O�ʦ*��biqe��N*���G�����<E������Ð	SJW+<�������;�v�q���d>����U���&��)�x���ep�M�c�G�F$<������~����}Md�_�J8ʳ���^rG�]�[���r��+�<n8�������Z㛦�����l��F��v�g�<0�����b��o�,�|����T��׹�y��T��'v�����=V[W'�Q�3d���MֲX�./�sɪ�����J�T�!��!���g��ziK)�kP�⹟e��̆4ųQ�6��D�ؘ�������FΥN {�~�6� ��W1v��Zxt�俑2�v\�\0ۻ�*��o_ cᗃ��c(������j%q$xڳ\/.�"�B%�	e�)�E�����G5q�h@g��7c�B�:�w���α�1��!���r�GҀ�(�����%��mخ&x�:!�9�ɂ��fӎ�g��\(���#��w����@�Z�(9&�vv�y���zFȾ�W�J�x�\�.t/i���}R�E�/�7�%��L��_�΢CG>�_��t�*WҢA�˭_�r��S?i�s���=�PѝP!o���B�X�:����3��V��4�"˗Q��� l:¸oK��S�z��3���C��^���z��~�y����{f-Vq8�]��u[�q����m��>�f��(�b���xNTS#aگ�ȕڪ~o��*�*��yu�m���uҧi-o��=]'�<��ި$F�,��ϲ��3L����4��Cߘf��n��͓ܯr"ݟ��&R�����h��t�D��)1K�M��j�ϷwO	i�J-D�%a����ݱL=�s�ñx�����:p�9A��ET	��7"�^|�H�7�7�O�Ks�	�Ĩ�v��8O�Έ9|�2v�nb��H(:�x����DF�����㼵��qyy�ͤU��2�J�`~���V?�+�8�D���Sµ��u��Ӷ����rX������|�N�A�c�>�i�.9�2��+f6�s.�����{�L|�U`��v�O� z_�$�"^�������P��/�XN�g�>�(\�ُ��v���p��BS+���,Ԫ�ADm�{.ZF����^O6ZUͪUlEڻb��e�T*/w_\��WI~��N���1 dgm=�_JLRʯ9j�m{o0�����`Z�s�\Y�H9�໧� ���l�\7/�4�D�7i��;����ְ���^z�yG-{���q�J��d��>�P6�G�L��Sowk�W�K�$c�R%�_F"&;'��"����c���&%P�
Fz�U�o���U��o��Jh$�@;�c��b�Vɘ,2.�m=��g�}��1Ӱ�Q{��e�����ﺂ
K��4�m��^|1FIW�guG�;+
��2�\��<��wh�)��j�8�!�hx��,ߡ��t�G��4�v}�+���8���+��c��ܝU>�;/��d��B� nx�D��L�3f��ÈofA�q��
Ì��6�X|l">��f��_"��(���j�c��
T��%L_(�?�	d�m�ֆ�t�2���I�Y+%�o�h��y�7}��|�;����z[TJ5'?˯O��=M�G��GrFj�f>�f-��m���$���1G�������
%��5�8@t߫��s0��kq�ۡ҅��-p���F�[�7�f�³@�ё�@���8gw�P,��u�Ѯ0��b߾hY�1Mh�4�]��q�Ta�S�"�������)̂���j�q����1eA���x62��rvQ�0�`�����^�r9�3��`֖��`��j����j�E`-%�(��23�[��WL��T&�+7�H��%���W���)�p��$��2_c��̝�ǅb��FY���ҴH潲�R�2onL�l|_�jf���Ĩ��p����S�3a�4N�be��	� C^�ٔd�!x�+�4��J���L����\�M�v�3�:"�[���`�o{Jʯ�E+��W��p��e)q�0�b�,�xyF�ds�˻b,�X����T����2�������d\��)�;ϒ~�BvYr��Pg�0g���[�,��?hc5U�v/7�k1P�������EK%��Q����GM�r��LJq��
P�o�\ (���V+^O�4�� �X���T2D����`�)�L�1������ۜ�;�/d�k��+룔���s$1����F�?ߌy<E_/����şԎwq�b��9L=R&��Z5;5���bx4�յo+1෽cbP���//g���*�bm'�DD�}�3���`ࢲ��"|����'R��a&hг@t���O���vw89������y}��js�Eo�!��kw��Kmn�.�ˈo�G|듩�4�0�Ŏ�#��NY�ڨ��Ie��}�A�w@i�/Cm%z��؅���y!�zGu��/�|=�j�uNh\�~�ж��.!�=�W�&��EķfȰUÀ�piL������m�ᱬ�����?& �ֿkV=S�"�=� ���O�ʄ�d��!�<�1�N�e�l��w�_�l���z��I-��$�$ܬ���CWsΥh�"n�t�z�Pl�ex/�.�$��x�+*�f�C7���w��F����ډ�+q�=*g��_/VM�z�y��\���L��k�B�C���E��o��	.�������j�f����+\Ɣ��6й)�Wq����I�a��6�����?�������t�oo�&b������5�N�gM{|��xl�!�5/��f�ᨗa�#���t�ϓ�`�c����}��|ʇ0��QH��9a�C�%�z����nq��E�1�t]�����␉�ʇ��D���~���Gd�q9gd�>ϕ���>���nzu�p��z���$Tl�ŝ�g3���� F7�۷{:��P�F#٩v�$Ve�����i��I>�cXf�=�#���!0+����z���+6PM���ˬ�=���_K�k����nMU�>���,�;k2!�w���6�v�_�j%p�=�9n���C���E��>G�ٷ#�mWD_A��P�Ҹ
�s��1��s��ǳ+!G��-6�,ᮔ�����;��p=�[鷂�X���BV��W���=���R�.L�7q�v��43�\�n���W���%K�� 8�ͥ뒵��^T�PI9�Ѧ�$��7������4{X�V���:�Țq�} �r����}u��yq�=�l�FN�����T<��JҵZc}`�r�Z������{�-���+�O����0h�T�kB����������
��]E�f��Q�Q���Zᓶ�_ܳ`���y��S�8��`��XkU�1v����e��&�����_���n�Y�֚ ���r����BG(g{8���"����t0��	����4 C,�B�oOianb �~LG�̘~� 9��t�O<Y��F�^ryq�Y��RS����`t�f�m���0]��-1XB^�-�\������^gt�1�l�_��E��x=
��z�{��1���?��WT`�q��=�3�! �-7;g�v�~}�P���r>ېWs;���?&�Q�q����qo�!Z�ڜ3[= $�w"B.!������[+�@��2�!S����g�$@� �lѾ��]}��
�W��K9}sn4 ����lU�-#WcX�*��w(�c�\\�9�+��\� �wn%��0��e�UTW�����	����|4�m���s��4�G�
�96;K�~�R<��*<�#�ƙ�3���C��˓�ⳍE����sӭ.�0��_��ng�h��C�S/��@��x`�_���ف &�����ÿa^Mm��T�cв�����y�e�L-�tq~�y��f��Q��~��Dl�[+ (c���:]��ڄt��C����mb����L�{�����O��������]���{�r��v�/��ߞ�w\�;�v#��P+O��[8�~�R��db��I��!��T	����=�+Fj���c=/!���fʩ23Z[�(��,��!�I��:6$�Y��㥺���� H�*f���M��) 3���g15�ؼ{���n�m�����&��8Ϗ�/\;q�/�9�R��CT��<͆�*y��J�^�%x�xЧ�|ԍV�/<6�`j*�|WY�'&�ɶ��@q�l|R��{�](H��C��Vbt�\�ڡXU(���APE@�s
��$��	J�����{[��C�Jo�]�
���:))"�(�\�7LYr��7�2�~"�{z�i�	���{��S\N�&�
�vlѫ�	?|�{7�Aό�����r�.�U���u/� ؾL�.�q����}'%����gzD%��:�W���d��܃��H�����OBK����q���o8��!s�'I�M���?�k<����~�6Z��jܟF3FpO\��x�2���u�D�TV�0-e�g���=8�l�n��la�}[ؾ��%2����c\^K����dE�\b"��6eM2���J�)�7�$H�O���ԣ��$�,�o"b��^����bƑ�r���Iz?�dE1�;��)�����X)DA��*x&��S��1q�O1源ۦ>쒜�J]��D��M"�IG�N�ru�]��'�E��<:.�]͈�}��7>�G�}풕� �An�R�Ӈ1M~�]�¹��z~��
���L
r�)ҙ"/�o�*��%��l6��ۺ�\�U�S��D���X���Vc�B�M���Z���G����j�J͝|жӖ�D��A6/A5Px�\\Y��)bx'�|�	)x[�^a��ݛ�!�u\���N�LٰQ�B͎E�7�h���Y���)?�_��T�ss�$7�ry�B��|�]���jT���z�o%�O�;\��)V��U*�l�7��*ɏ�ߛ��룍���ٽ�� �=��!Ke�	�с�0�4�����m�{فrE���1d�s>�
��3�O��;�Aˡ��<�L.ll'MN�(�I�Z@����̗֋����5:"E������B��V+Ǹ:j��KHp��=}��bZ����ĳp{2�u3ٟ���w�%zQ�	�#�-�Bo�x�d%�M�b�n�Á���e�,��2�I�&�_}�c+�,��1��;9�%�J��5����\D����o9yf��9���?�H��a��]�@&��z�M�ZeRQ���Ј0n���z�6.��m�|A�e��m��q����0Sfxɇ)|���k/\c��6�S��F��`L��ι�L��8� Բ�Dlo�N�ɷ���s��ӥt�?���}�fp�_�0k(T�?ũ,P���#e�0��`��\������Vt�l }�z��*�Y����!n�|9��� }ǟ�L���H}��r����	~{!κ���̈�C�Ymx����@
�/c܇�K�/��E�1�^�n ��wh��!d�O�����~��s&3��%�RY��QY	�1�f�����o*�G˝1[ޗR��s���+7!���T�TPX^����o�H�h/����ظv��.5M�Ҹ����X�4�@g���t��`�����* ��� �ڧT3=v�
�`��	����D-K��oo�(�W�$���،��l���F�nZ�V�'��!��n}]]�K�L t�ڏ�0�f�XYD(��R5��*o��p��?Y�P�����p��>��z�jq�������y�[~.�,����8�WA��%t{/<��R����E2����.n�U���W!#?\����t���+�qbF2���>���ܶ�ȅ%��'<�z��XqѴ��5T�)Bx��'�/��E��V`_�nqd[V�f�ӭs9�w$��D��[hӏ���ŲEnp	ꠂH|���o��32Rd+k�n��,ϗ�m�O𸘍��!Ԯ�h����%���{��*��n	~���y���ǜ���f�A7��"��}�H��]Tþ)��i�c���(J9^WR{�E�B���|�WKy:�1n�d�=��lb��㛫��
Ω�~����Ғ�������ʹ�@�}�>-iVr8�'%�<5��j�����MqH��
�:d���)q��=^�0��ũ��Su�hGGLk�K�1����/XO�AhE#Nɡ�p�Cv�׆�v��+=�,�}k_��)��=���re�fir�J�L:v�59?��C�H�bw���� 6>r���ixN�����w�l��q^��.�&�=r�Ly���wis��`�9ZꏱO,���.^���<��l{[�y�����,#�u'���yP3�'}����Y⩙J�,�B$j�=������%�7�{*M�8�ɵ)Uu��Ko�C*ֆ0��J�*��� )�'���^J{��Es{��R�gO�e�{�L��֒�[�L��
oS������	gu"aԋ�}�Z,y��d^<6��+G�Y��`rE+1�:���іr#$��o]B�L��3�B-�j:ʗ��L��u��ᕫL�s`}�1��\���V�-��6�����[��Soh#M����OxȲ����^��i�.��a�BD����@ߒ`��2E��:z�&ΑJ�ӗ��H���R� �5�	`+�<i�,��N<M�a�
�4 ����8�yD��k��rЇ ��F=��l�ȴ|�!����8B�c���߃�R�G�R��Q���ְKq�����o��M�������t�y��G^K�.�qW��h87�l��:���h-7<^�*���:@4g�� �e�k���m����8�E����u#�sa����ʰ��oMJ�X�@��^��{��.Ŋ;��^���J���+H��+N	�	��������~����df�9�cuX�kI*��N.�c{Q�j{>�����]˖UJ3�Z��@�N
̿ANԘ���(�c�1�Q�T:��j+%@�)ߤ@!�2�b�נ�
!��.3�V��ɦ��3�S�B��r��3��݌�_p�wV�o2�*�4<I�hm��^?�akYO�hBƠ}I}ǩ��K��k�w]3�������,	��w��Q,C ���������Xo�t�E�Ö����qƅ�Qd2��z��9R�b�mWg<<����;�(v�:�31z�>e�"#v�q���l��ni�lT iCw�gߑ�S�9e��z��*@`#���,/+G����@�=u�Q� � ���I�&��3Z���԰x�n���%$H��c(>�|#�ԣTo�͒-�b�	���$�:�����IIU�W��w]����<�N�͟U�KH4�H�U�M��\��6t�9]�OflD�%}�`oE��E$	�o����K�S�=H�%��MF�_:���O
�����d�LFD�������/����۱�/�r@��U��y�pY<a���]��Ż�B�J��)b��sW�?s��*O�J�3��ˎ��S��TI��$�������z�Q)��'�;H�!�U��Oц�>^���j��ݹi#|K29�d�{�>���	��S��
���MK�&<˵C&���
�� #,1�>T�8�S����}"D6��-�����86�r��Z����B����f^L.�JJ��6	�ߞ�(�uGz�����N��#4.�Q�+.�w�,��] �ϐ�2�������nר�C��_u�V����ICA�k)?��>�~����My�e�&�߰&���UkA�A����Ό'�{&HY����<t�����F񬟞-�lQ�%��GN;l�*�F\�\�8��ɏ��ssǂI���5����s9�����T%�Ee�j��4�1����{���$#u(�<o�-M�	1��D������L-�K���cJ�.�.�ǉ���?���<h8͐Z������s�G�Oi�����I4��8�z T���K�&|���9��;S���!;/u��E3�mo)G�kԥd���Cpe�f�A}�ɛi C�v�)���m?�"�qV�/���o9��/�Y6��X�o����RdE�5���, �4&��V"�+��r�����?��DW���g ҟ�[�H����6�uˇS�XJ׆�s	*���P���hD��a�H��Ml����2�+��b�MB�5i�ߏ�j	�%��F7��ߟ��J�q���7�J���X���'ټ#�e*�t�(�­Kb�n%��������&OM��!?S������֓!��u�UUU�d���1�Ry**O�[>n_���f��S��v����YZN��M��z4'K�Y�}H�E�;�A��(HcP��7�?xK3��V�� ���н������c͏�k3XZ/�Y�c�v�E����#XF��,Sz��+rږ������FMO�H�dI"yG%O���i��	HA�x3a�S,L�f�
�'w:C&��UQ��M(�h ���p1�ׄ���]U;������o��X��YA+���Aw�,,H8��c�~v���������.�F1z�+�p̘�Z�/kd�S��~o2��(c|(���!o�s�{��!�,+qn�>�[�ꪀ��+�7jZ`�jD���j�3�c4!��a�7Ϟcd<`!�k1J#���o��ow��淿BzC���n*Cι/k�w�)C.�C��<�3$p�u�r�P��¸��ǽ���ztE�6�5�b��`�l�i@VZ�bk�hJO���n�@!�k��A0�/JZ�1"��~�����"��w�T�r��kB'�x�A&�ߴ��=/��՝��3���^}�b���z3c����[� ��fES�#ǭ � ��CT�ڵE?O4�k?ֶ��.�9O6���t�]�}��z'�pQ�N�*�][�L�72IV �n�����w�Nԋ'q��$E���i����_�\�h�P#���+lV�hl1]iD���,���_���X�~r���ن܉<��@.O��Z�[����n���"o�>�ӄ���Š\�|f~;h r'����1Z�VH�"w��n�
^��P�*	��YEpk^%��`ҽ��``]���	6TW��U���^� ���^*�c�Tۚ�RTE����a%"�I�7~�פ%���N��Rj��M$� č�&�o*l�n��
�� 5
,ۆ��Zʼϵ/ģ��0���y�����Xk���b!��qc�Nen���]I~�D�V1I-. � Y�>b�lT~n�yr���ɖkˀ��X�f�:�1��K��r��B�6�:�$w�s}@E�J;̵e#^���G5�_��kH�7���M3f�s���V8���냰bBb)�O��>쀌a�vq妵���L��8�h�����F���ͮ:�e/�Q�Q�����c��w'�S��i� ��p���� ~>4�$'u����^7ffm]xk�]����ψ�<��Ć	{��1�0�/d�Ҳ�%�}"��̳�N����:;��/QRY��yӢ����T��b>��͖쯜VU�G�a=���Z�Ǖհ^u�QJ�ņ*�L2D+�~�4�%���n�/���y&������j|�z��l��s��Bˑ/~��RBPHP�}-�;��GĆ�����Ge�j�C{����+��I�+���>�9�X�'tt��:ݭ&�ǘX2􄖴�DE*a��^߇y����XҬ�aB�
6:��lZLp��S�����.`��M%���g���	`��qi�W�A�E�&��>S�zMɋ��e�����Nڡk�=kJ��s\�RXi1 eY�][���)ET8B��wgT�X��^/�u?{���c��l��;	G�JC��<ⵚ�A�6�m()�9�\B����L��=��ս��u��M�vR��"�a����.i��<���u�i@���Q��
6�R&)9��x��2�����{5�^g/���8���y�5niC<���0X�'����P[;~󩨅�gkH1&��B	�o`ҩ�?�l�"A���}��_K�axE���:��C��7ҡ����$������⇬��w�2�%I�$�8Vr�����>���w:��$咷���@٧��W�qA���2�0	c ��;9�y��.¬��#H�I��D��(��#�F�/����s�,v���-Y��D[C���U�ȜH�p-K\ю&4���_����S\^�$5+��^�P�a�����߮�$��~�B���Ĕ�5a"*c��C�2"˓4�_�2��}�疉K"~Ƀ	�bˋj�nd�"����R�������:�������6
r]�?1��-]Ȗ�.���`��8����-��2�v
�TT#���V=ڍ�w�K��]�����]�c� r!�SXV�}ƭȥ0�`�="��/ 87t���%ñ+I��ЙL��ޯ�����F����Z\{���K�T�y���P�T�%���F�x���9i�+\�������5W���mۣ%Ҵ^�N�^�2��`���5L����k_����v�����a�1�3��N�����V# d����inF|�^��gV}LE����ë,n���vm��
?�݈���hV�%���`�E�y&���g�Ȓ�u�z��^Z6�L~��䠻 ����Y����+��V74w)(�e��p(�+�E0~����hu��c%���5�im��ϧ^��U��δ��S�.�ء��nvЮßȯΉ{�N��i~,��j��=�n�/�S��]�5�� ��ݶ�DA�VW�*�i&����-�ݧ��\������Е�"Y��a�\"-�NJ%�����{�1{5K'�2�v�N/��m�L�!�B�/VL#(Ƈ���nB^�~5g�y�`�+�٥9��LF��mb�|����+(�i��S�����`�V�{�(I���H�,ט`t�5��hh�@.����'VW�}�jR�4˹9���O�=�b��� ~��7a��l��<th��t?�c*j�F�H}O1ޝ�����,w~E F�|��E�	��N�G���ͯײ����[h'��u���3t�go�Ǽ�r�^���L�*�<�.��wNx�D���rա<=���(�X��f��̭�+Sfs}~TcMNZ.�ȗ���b�� ���6Q&�":����k�*����-��kvC,v���-��3їI�"�	?l���Q�z�Y�A4�W]�����a�q&��=��4�ė�_3��-���|�o�� ��O��Sr.
�Ͻ�éo]5Lݏ��h�B5��[}�-���bYۄ��w��i�z���=Ř~t
�[ޘ@���풴�W�`���%{^s��o�\2��\�J���=Qh����JN�:���@<UD�+���[��X=�k�8����rt�K`&�x�nd�a���QJ�$�?�
j�u��5������J��`�)䤘�>Fh90�1�Z��+�J�[��;kQȑ:`����ί뤴v́o$	�J�mni��_�<X�ȱ�I��C?u�zz���C���}�Myc��#T��������y�yĝa���T�}��0�3��%�%ޭ:�I��!x�4~�%/���c�в�vS��W5'�>!��Z۽05��J�uE=d1S][�j�ק*t��%����LUJ\�`dDľ]'����zi\=2�[�J:6��H�ڰL�cU�u�\��x�jby����U�T�w>%+�8�0�_ċ}{@R�ݘȣ�+���~�t^�;���Tk:�b���K����/2��5��k}�m�V	�髇?Y������ 6e^^Ϭ��?���(􂂼�=C1�/ec|f��+�=�'l���%膾�sp4�c��>�Ƶ��Nה,'����a�wn�I}��R������=��y-�}m`M�?u���E@@�b�Ď?*�td�X�"�m�� �꒭5HL�O����/>���q��y�I�t,:~�Cw�+vt���qSo@y΃�v�ow�s^��QTѕ*�V�/)'�Ε�e�Q��8~@0j��M��� 2V�>a�b��.�{��cV���{�>_<�bw�rr�v�췷8hC�(\X�p�- ox*��U��UF���_t}{Q*P�z������q��C� �EG�Ԫ_=�wy���~8nH�KK{~tSm�c�a����xir����������d֝o�}����(�Y1ъi��8��-H��sKÏ���~���D�E,.���~!�6�`�_L�n�@an;R}L�%5��I��{�h��8����t��戩F'LX4���E�ޟ�����v���N�DK䦼,ѣ �uw�:��멳�PV|=���aINRL@��5q��`(*[��<�f��ӺSȰ����QL1�DE�}��Pt����+W#�������V�Q�;B�'���x�Q�����B~ ow�����!��%t\,�vŚ ����D��ՌEm^Y&��~{�o[S�,F��|kc�:^�Ы�#w&�'c[R��)�jݶoU:.��̵�p{Wra��J61�K��B��3�¡
�(`f�
L��_����J��El��oG�}P�����^��K�}Ô&_�Beպ�G^���R���1��K�b 25�
��aU @VM95œ�P&�UzC������0�����>0���	��i��sr
����թ,ҋk�?eO,��4O�(� ��~�y
���7D���ŚnTR��F�勵�z�R�r��u^,�	S�O�\�t(R���oxZ�7�1PRRb�����f�=�{ۍu��~�����+F�	���ah�}�-�V���%�%����U?��,N�����j�E r���}�Y;������g�:�K���A�Ng�������|�� &Ԫ�^��&�����X�W��L0�	�,���ﭘ"����R�u6�*�H���ȇ��9�vxeh��ѵq'4��}s��Ӟ�S�s��V���1�a�髥�Ӄ?s��|c=@�o�y���VCSӰ�xY���s��9�E���E���ޜR�JF!��*#��l�����z\&�Y�����g�?�*6q�A�*��hZrumX	�}�u�)���/'���}�"�D�;��F�W��D�A	�*.א7{p)�����fb^̹?_�d%Y̵��}7
��	Vǥ^�,gU��6��Q�t��*X��gd�w.*����lI��9x�w��R�jV����9%l�����sU�=�X�2T�y ���V�^���.�
Sf1*JЉ��w�Dʌ�I�i#��n�y����vk'3dB۬}>�r��.[J<X�ӝ��1ɗB6H��߷��_�r�`�^B���4�_���M�����X���}��������L[�y���t-H����m>�c��db�c�}�S�^[�,�sƶ��;�"~�]>����aD?/�g�ϬS)�f5Tb+^�v1bz�����>lϟۖ)�rz�A�5���9/���� ��ߏ9/��G?4��O}�\�6H���Bv,iˀ��qT�5N0��8u]KK����X��.�<�v�&й䓨����	���d�����Ŝ��UPP~S������y�=�"�w,��脈ݐ��!��%�$kJ��cs�����S�q�;^*��)Y��x���<BW�\�A�[�s�teUuu}W�v&��4�r�w�'���sh�?�<��	d�s�6NNy���D�^�B���q�
s�B��R�������S�|Eu�x���7y23�hb�]�sq'gdx ��h��3�(��Xڰ�4�}��e©�}F�m��î�1�I�?�.v��}��zy'���<�O�P��Ӯ�����j��]�OT�U���T�s����7�Yæ������_?T��g-; �P�7�����S�ªāb��{`�Z3�ʢE�il9�j��	�r*��gP��i��&���.RB���5�G�^k#*g�5��#A�i7��w�^ܒ���!_WW��w�TgB��H�%����vXX�ȷ����ܭ�23���M����0iX%p6������Z�x{�%3'�Eӭ�$�팱�U�����pHL-(2�j�g�\��Z�]N`��s��C�˧JS^Ïٯ�]���NE�{'v	:��H�H���>�Df7�uq�m9;������G�(����n:Om׵h2x�};s���z@��/�9^�����}�r����-��]u��="��SB�]�r[$wF��Y�>��-�",[Tu�I��������23���FR����;e�V%��/�-��e�E;���7��j�ղ�T)V/+��r�컦8�_k�l���3���UtL �A]�o�f�Ѓ�~JR^����+lē��*��^;]me'�)L��,hϳ�[F�;�jk30K����/�a�_������S0�����B	�b�U�'��%�9~p��v_��PU�IuB�;)�`(Rѓ������jZ�����Pڀ�����R,�{Ia7������E�hFa�'E!j�Ev��1�WD�z�����_��W�Wi.車!���rgWWو2=�As�r�����i��b���hl߾BZY�,���5��ʡ[.�t8m�z�#c�,���#{���lz����j��th�ϯ)P�0)���P@Ϋ�`D^�Np~���ޗV�/��-d�f�ƍ�[� j�̙�f�2o-'��'
�w�h;
F3�zz�=Q)	�,j����B���S�����π,�ǔ���1�����z�n�f���4W3UͲx��)���b�8�l�3���{�0\�6��K�;˘[VV05��rK�T7n�z��U�����r*���3Ǵ�H�T)�L(�3�˂&�AQPH�&8���e���᜖i����	b�ݩPȩп����w$ݗs�G/G�5$�Y����|P|Q�*��Q�X�8W1��J*&������ Z�T]FFs����vk�k�I{���.����眷܀-�U���;�)]��l a�[+�!;[GU��f�!'�k���)\Ɲ���è^��Ӹ^�CU��k�G��s����MR��C����bV}:������	�uSt ,i5O�m@��?�ZG�7@�#�ڭQ��Vȥ�U�R��)+|�L��#Ui�u�ܲ�(�S+�U�tN�1;�Z�{5=�hCc�*��iy@�G���C���9C�����G������仭d��D�"�Y�t�����M�zr�2���:fݢ�\W��d�Ȯo1���1H�6Ŏ+�X6��Q�{���qL͍��^�����Q�qM��O���������ͽ;��"�I[>���k��_�����?�R�璖p��	�ƪ]o쵔�=�i<��-��=���D[-$K�7��%* rfe�v��O#�\E�4�M��~�H���g�bW��5�XSS���u�WOC��,%���P�a�WC�2����V�H4�-Z��a�u����碠�s���C0;;���%\��h�]P|��n�f�ϒ�S@�k˯����]��q�jD��;��MN����+�w�ᓩOi(��iv�oa�%r�R�DXN��7�鹩[5m*I��D�++I��Q���ν�A�F�WZ:Yc��\���ƙ�P�|�f� ���,��jX����ɕ3ݍ�d���bӨHb�)�!h�� 0Tc6���D�J�6*�>�z�G�s�M#@��������x�����$�0O]fڏ9�<�H+�a��#�H���=�:����z9�׃%�Ǫ��?h�_��<��I���\�q}�P �D{�y�{_�O�Gޘ�'>8ڢy���m�B��7���?���X�_(,4:�c$��ϵ�R����M���)�r�{O���A��%oc/�#Yq���o�N���|����P��M�
�+oj���O�Q�46����?����[^��ܤ�p��*�������V;�2����g�����,X��V���	���x����Lq�%L�Gp&F���
�Kg���9�rvu>��	����O�Tم �#�x�ŷ,�ǯ�Y��e��I Bi�yGn��;$<�1(���xt�;��fG~:Ug"i� �\�$a!�t��2j����uS���t�6�
�v,�βf�2e�^��,���%\�����_�~�՚���d؇q,j}4\#��n���њ��}ۤX��w�8����X*�`=/Ϥ=�)<�<S� !|�r��|�x�xw���h�qt} +)ܳ�>��_L��r~���A�{A-$~��#*X:F:�))M�:-
��yמ��;jr�e/��u_+���ta����5��G�#�qay�SzD0��r�K�a;3�����e�/�;^��\$ �85�voY
������A�SI�=ae�Z,�f���� #zPI���V|��1��ޒw�l��Ud�k�C�ӏo��	D��R4�To��ܪ�����ۊ9�z�1��T@3��6Z�w6@"]G���V������zrw�`��u!�7�6���~��g3�K['�5�^����P�Q��v��i����=}��U1��mSW����FgNpx�B��nZ\��[�ܟs��4�EUB$
�]+4����YH��tD������p B|��i������̌��٤3�X�:��={8+�X:�L�:���Rum(���ũ�8�/bl49����ҋ������jk5g`�c���Ǐ��拧�v�9/�`�����q���D�G)-�FŲொ�]���w��	e>b�/�^w�.���}qdA��C�EUw������uA�@~���{�_2���Fz���;��R�B&��Ы$��%�A��:U��y<�M?�}L��tS�#�A-5r������\��l4ys�\�m=�!�D�G�4n�}jQ?L;N�_/�����(��Ԟ��u)j�����fj��L�n���|�_��C}4X1���z �Y��"�Wյ�����}�<�>-�ӵK���y��Rǀ��lǳ8��� ��!�h��ܴ�:`�fN�%�H��h��7����i�����w��qt��&����eh+�񯓨l�@�+F�N.z�/a��}%*�a�E5������=z���сXU��q,�z~�����i������<Jr77����7N(�d"���w�� 6�@��1��{���Oƣ?����,�M��8���T�Q}��}��Q��!�������Fqc�"��r͕��O��?�r�Ё����ߠ容����b.�y�[��Ҟ�~�G��#�����"~X񖓾���x������Xa�\Ѡ�����2���������bT������?����S����4w��̝0����o���pֿQ�>)����i9�"�S���A���hI�8&dxr'ǡ�ye�鴈�
�_S����c3 .��Ŧ���T���F�No>���o����������>��7'����x�$���3��&?���3�*;��}��-����l:t�#�(�|�L	Bɰ�d�� I*X/�=��h�h���!�<���E��O�:%wNPbx V��'!HJl������DB�%1�cj�og�MO�|�<�<�T���QK�8Z��,�+0V���-��r����DJρ a*P��]_\,��V�2��[�PiL�{�%�F�F֠d�6@N�"L�£�#p�X��dİ�U7KK��[�Z22���Я�y1��$PӲ�0j�f��>���cx�'���I1�Y���j�nwt ���q6&�)f,�6"AT�o��w'��e��K"6�����AلTfƝSU������Z�2<ۨ�{,��#J�e�P^P�N�c�5��ҧ�<��!"�i��-G6��D�Hw��#�i�������i��c@ٸb%-x��@Ic4���u�r����)(Fk���Q�D�W{M :GxKe��T�-V�Zpe�8 �4Cڲ�"�ȼ�2(�3i�����FM������Gp�z��[N�'	R����*�h�*1�a�J��'p��RԘ�7�(v��a��/���-MvCt�Y;Vzt�#wXdA ���k5�q�t%|�z��MwBm��*�R�J��xb������sy������"̃7�[�*������Uw���Z#j�Zϊ��BZ�Y�kV��k^N���Ԍ��-�(�l��r�х��G��uk�-Y���J�zP�PS �=����f��B�:()j��|�?q akTz�)Ô�a8��������dc�)Lc���#�q��l���h�B�玅�����l^�Xk��^���u�!�;wH����f*G{�n{�7h28�.���c�H��o^�Rӈ�}���A])raږ���-շQϋ��Tk�ޫ6�ӄ�I2 #�2�Ӡ��%h
��rP��6&Z�h}�N�r�_�I���d���`3^�����Hۦ-Vy���b��\̺i�0��th�����X�|� I,���i��G����~n!KvhR����
^���+���B��`d5��(�^��)~@z-��ȁ����U�ylфL���ۙ�hlioy�7i~h(�T�B�1����k�|��
�2)@ɬ%6�}��p�>�����&��җ�奧�ƞ���*_�4l�q�W��xj[�^,=�}���=���0>d����o�����ot�A{�Dg�M��K�(��s�K�[@�s�{v&U{��d������JR���Y���K�ْ�bȻfQ�b��Զwɵ����D.j�O�Z�(��32�G��/��'Ey��责�]d�~�i�m[#���l?�ܤ(y���c�����z�W�m_����@��(((� ���|#	��\���x��z: ����WL�~�2��!q�Xy��%V�6�����oC�1�<����>����ݣ9����ю�vf����j��0��h��D��dC��{Jr��b<~�|*����_g��|X6��CA�p� �R�0&�����u�����R���Q{Ҋ����7��1�E����Y���@W����CEa�'��$j3з�̢ޘ�֩�}�����u߳|u���>�MF�i��(9��O��������"�c�����q�_q�`�4��6Z���� "�����=`�o.']RȪ��I�SR��'��-H0���Z�z���:���A�ᒯ^��b�c�f�Ȑ�L�����.�E�/��{'��<�X���V�ύ��|��f�Qn4F��U\�^�����a;U�3�>�����������@D/�6�1���?c"
� ��׮�{�RW���;S{�x�������C��:��HFQ�:8��%�����U��X��ء��;QM�����������W䲯�� ���C?�ػ����ȁ��nX�AUA����0��l�=5�D���`���'��B�����w�Gm"S(A����osʇ0F��w�_%RQ���堌}1D
Xt��o�hܿo�.�X��v�F�~	|�hڪ��xᭇG8���ؽ�s��8����y�\ss��s���5D��Iwp���;��k���>kq���&]e':��H�����������4�2�hT�O���/FH=E�()���~i|�}V�}9�v§�V`I���A��`Hf0(�YJ&(� �a� ��mw��f�K_f��\WCo�BK��>�L��b�8!�Av
�����A�׼Ԉnk�r���e�MF�|8�h��e1�� W�vy=��`��n���z�>Ƶ�H�J>�i��7ѳ�/>N4/�L+G"b�g7EM��ʣ�����ۗH���dA��\V���򴻙�Q�"�)��@Q5���b�q)�U����`�Op�����68w�z@� ����o��3}�@KHm�W�ä�2��P!'	Q�R��;��n�~Fy���P�G����t��c���m�[�b8r�r~ر��Q泷Z,Y�M"��ua�ZO~��XIO�bϣ�l��︁������x����K�O�۳��9��x,X9w[wz	�m02=�� ��b���������H���Ő���y{�јx��Z���2>;JS��)�D���o��Ќ�r`�i���o��W�V���T֞�v}���5��~kF��;&�$_�0NB=P�G�BWTz]��ʜy�/�s��:�~r����K�3_=�A�Z��r��!OyF����*l�(�y*4�跈"�&4Hm�n�k�p���ހ���� ���F��!@�SVx���3,�,	��ܦa�����W�!�4W4w���35fvN��
�i��8����a��wi���d�Jt �����`�����_�s)�?Sk��в;�Ӂ�w�@=�K���im�)�_���x��bYa����mj�R�z���*��m���z*�����to�#��I6,���������݅��ww��<'D��Ur��]rz49ͼ��G�ʅե�w�l{,�1��?�>�9���]�<$D��v���gGD�TmB�:�5���p� J%B �N���O�{�/���S�4������Y��y�	���
PN˲��0�`ڃT�d�D���	�J��hH�kH�C�s��u�����B/Е�=��&ێCt<��ڪJq���\��1��=�%Q�n���Z|/߯.�t�#�M�<svj�:۫U;�<w�'KðW/���Mp/��'�_3���{��rB�,�e�)C�e��v� �-�"�M߬�1����G3���.�~�����}���B q>��O��_�N�H��׆W��etS�6&�`$S���"�`�{� ߜ����$�:5|/.�s@U�[I��D�+��C�Ԕ���et��	�P����~ݧ䌪�yK�"4��Y�g���[��y �����W;Y�y|�w��d$*.�#q:.:����e{�!b��9i"�c���+���<�f��t�dr.`p+P�I>Q�J.�yA�!O�<�3�J�Y���J�(	}UtTP���9��_�6�'����)Q=��6^��2<s����:�_����~�h�{���U �4c�i`~�j�{�gv��
,⑻�V��R᝺'����܄��Td�p�(�<�!H�HxP���k����h�Pr��e�y���"uב.��.�� ��暲=�u�Xv�ah�]�Z��H_�T�:+e~�1*u�J/���W�-h��1'�\�C�C�����s�n���,v	1�x�fپ3믰�j.��d�������岻���ؿb�����+$MM<���E�4Ǚ����=i��?xPv��g�u�u �b�X�_]TU-,ϴطOi�1�n�^�GfH��^�a�bЈ���J�uf,��O�M ������4ٳh_\���W�>��)8�6Fkn�E������o�߆z\e��ϱ�Ĕ���T�Cv�|׽�w+���߭�{l>�x����Ĵ��?�uQ]<�0.F�D��&l�`�Z�V<i����o��]�<��S@ dxѺ�q���!c�`��Ȅ/���0}�';�Ng�!WCv�k]C��u���S��i��<q�fR�H����IW�fx��"X�_س���`S�T��{��sk���;"��cTrt ����꟣�:a@�ص�*N��X�Z��t��x�%6aZ,������М�AjO�p���\_/�:;��Y�jTZ�&�D0N��#Ł������;��9�9��J"s�9���V��:^���^]Ji3�	�A���u�Y��#��-~W�>���)��ΞNUUu��^L���M�wg�P�,m�9�~$���$^�V]��#�k�j@5^�k=Qp�qb�L%�S��+,�Ym��tފu�8PxI�]|G_
�����qe����cA������=>3��C����^t�d�>HH󕛫r�_7�(�`Z�i��z=atnN���{_L��� �'82x�����omJG���_�?Y4K�{M�q��N����6U ���qFc�A�u ��{,F��y���l$?$�X.�t	}O�!�7�
�(alw_B����7P�S���m�#p!v%H��#�<Ե���5E���Q䛭$���X_ӝ��[�Wu�2 ʓ��V�`�:�^�9<#d��F����$c���96=
�bƦ������oLɜ�y{�+:��~Z��@o�'�Q��C����SX�T��#E�'Ȕ˴�gr���"[�Y���
��E�u(F��h�K����V�D-�z���<I�+����̿ʚ�*��4���w~�*��'�Й�:Z������44xe}w
�IO(nY>'L&�(�dܪ={�<�/]�~ӌ�����q/�H�ڗ�g��v�1
�9 ��إ�_*�~%��2�N�+kJ��bdUn{Ff�W6K�k�~3|O�D�UV*�f����ҧ�d�|���^(�R�O�~����;��]G"!w���x#�%S����\��}6���\.�N���_�=�ֿ���5���fL�BO��1Û^�H�	�߬e��?֕~�&�߈��C!�X!�|����	��f���9g'�]9�x�	�����ʶ�f�b�r�C�h�����H1�����9�]��4~
hu髮q�hh�p3\���X-)�J6}�ACD��������nӢ�2���۞���m�iI��-%ƞ[ޤ�A3��I�/���^����O�{��j]uKt7\���Kft��>*KK��;T���/�eY�'�x��b�a��qqw^l*?��E܋/�n썃�Q���g��Õ�����x�� -]'���f�o�n2G���P�M���膬�U�	b���κ6.�:.��o~��%�9�������ϣŦұ�4��^ӌ~�ƹ�Vh��cv � �]LA��y���,�lB/��[�1#y�h鱶dྒྷ�z���Dz���Ҫ�ޢ�����n�3���9qTd���I?�wa�&�����N�/��l�.�-d��v����VZs�F!ͬ�a���E�NQ�0ē�!�@{����G��g4"����n�ߖ��p��8�%�N �Yz�͚m��;�/��\�����ܲq��NBY��.�;�7SX&˕4�w\Q�D ��ю�Բ�� ���5y+GQ�l[*t6����O��&ߎו����r?����4��B�(�Z��o��"J�;~���ݽ�ߘ�nJ�܇7��z_�JL_ؚ�ύb�����q؉���O��b�J2��ʆ�
H�X׈S@���𗻻N�w����i���S�1��Ź	l��m6����&��~Ǳ{uoþ`Kl�p��8�����*��ҧr $�AE��ɪ��Č۫
�Q�,o�Ng�!����3�+�ޥT���h��H�ԩ�����ܬM�ڃi�k]�H�7tA&ޫ�g�S�@}Ʌ�Ǘ:S�<��tvJ��������I`����z��T�('z��&D��bD�\V�+�d�k͟urZ����0Z�y�?�f�)���k�F���}�T6�L�K\s�e�"6�=fa~�].��,RS�',��������1��)��k	=RQ:G�`e-S���@:������{8q��NSt�/N�'��k��B	�2�6����dr��	^x�3����|�8y�$�>s 6Q��S��h)*#}�*3M32ד��u�x�	^��gy饗x����]�Bcκ��%(KUA�SUbJ�GT�L�������:%�K����Ǘ�n8�'J�]�R�E#�F��n��{��~�%>��+��⋜8~�A�o��������%�Z�� ?Σ"�w�I���˜̯��hF���Jf�b6k���<�(��c�֏8������!%?�_�pID�G���±Q�\�y�ë���T��tZ��Ҵu;��'��X�ɩD[� �*ދ��St
J��8����E��D�".��M[�x��� \��C�<��.7�B��[����k��Ɨ��E>�����]���j1�3T��hV���[r�Ge�	H&e�*��Ah���b��R|T7���~�H���E)��h<fR�y������=����q��������h�fa��HP��l����y	c�F�P7N�>��>�
_��Wx�ŗp޳}�.{;��()�N�j��.bb��J��B9
�;�"(<�B������r�W�\�$ש�gS":�.�B� �<q�q�����w�wx���4ák��:.���w_����g���}f9��w}ՈA�H:����ޟ��q\��{D��B�����խ�����7կ�4�������%U�J�$��&n H��="����s,�3�	$J���ϐ�����ξ�Ҙ
c���\�_�kP6o�f*?u��{;&��d��e���p�����-J���4�@Y��t�p�5����%�tz{-:q�=���/��m5{`5�������W�� s�ȴ۽�,h�D5�6eM���U<�X^^eue���uVWWX^^cee���%V�V.�j��਼V�)��-.:�`���Y/h �L�*Q��~Nw�(��� 0m����[�մ�0p���yﭷy뭷�p�rL���i'��!'-d�K�P���lQ���4���P9�U�B=`qe���UV��8qb�'6X_[g!ԸAͰ��(�䝳����+�sD�J��DF�:x޸��/_��,�5�	��kd���SYO'Θ�$�$!�p��E^{�5�~�mN�yN5�e�B��b�浚vL�I�(����*�+�,-��T�UUQ��lT5aX��!UU[4.D_��Pŷd��v2����Ƅ��ɍU.]��k�]��ɓ/T� �{�fI��ϣ�����͌.y	:*����啝T�~4��g�`gE�w8	�z@U�:������������[ceu���%\��z2��<�=��̳�[Jh��o��l����Q�����/Li�Yɦ��
�|�8d��N�l�h>ER�"uH��B�}	��)��Z%5)&%��-�['��`�A5PB4���%NU����^�d�u0Ui��S�+M�3���۫y�J����43u��<�����Pf>>3! c�g&�YZ\����{���ENn�$��>BQs��jn���eQ���<������UU1�j�@������z8d!��2��UZ/7���!��"zg���Ꜩ��y�y��Y?q�j0@�Q�,e�[�c@=���$�R����.^��˗_��˯���@�+�-���nn@#@���P�j]�A�V[��lf�P����
W�0�r����\�����2�2����D.y�����+�{�'�ש�
�9v�i��?�ft��t�V�#k�.��{��Úvh�zʠV��S��ya!x,
�ư���z0`02�ԕͬ<Ma�e��u�}*�Ҍ����O�L��k�������
ۗ�������)�Xp@J�صSLJ���3Q�q�]�m#�H�9��c�.��#�O͡�\B�5U��Y�&�������G����B�
5�@���@��;J��k�����Y`���ڑ���p8��(�q��4����HB̑D���'�y�ŗ����q��)RJt�Ҧ~�Y�J�)%�S�>X��'��j���Mg��Rd��ÅZ���H>�u�.%@�V~�y��{Q�bu��_z�w�y��_8���"�	}8j=D�/��5�&u�ɓ������K�<}���i&��I�xfRԟ�YA2P��`8Ԣ�.(�^]��|��]��J�PQ���W�-!'IɺݯM�&)eq�0\�T�t���^�����/��P����t��	͓��CY��r�/c��_�k*0������u4���e�x�FN]*�qڊ�
N��J���2iMe�U���F��d[���G����`��1�`\����0�>�����(�y��؆/ı��m%�TG	��B��<2V)�f�`�qa@=��5��xW��5�I��3�C��4_S,�5UU#����/BE�$�f�	#��<���P4%��⥋\x���;��?M8א{�M��R�@p���Ӑ�iG���x��(���^�TI= M��5�!��!��"��A#�IMkx`��m%���'�	�O���W/s���Ҭ
�u}C�����}.����L�Å!gN�����\|�"+k�t�%'�]f�@��^�����',,0����@zn1]�r��a2�k��QU\PF+ޫ�*%u�f�u)���HG�j�_:�K/���Y\Z$T���y�?.<lu�14g߶9$�fg�$����j��������p@C�k�����\r��pD�z�b=Dj������L���t���(�{p�<��a+���'���gJ�H"������!�I��fxW�M��b7�n4_ID�\,��9-�WUn�XU�����kw�&�+�t-���D!3X^^����\8w�'֔�d�a�^�*�j�N�r��*��!P�
��B˔a�u�W`��D���#y��淆aP+�Ι��Y� ���'8�.f9���>���0F�7�e!���u,еH��L�Z]]���t��O���5�%j����<5^jC{�vU5���B,c�|�!L�Yѐ T^k��������F�GҴc�X���|��Y.\��ɓ'Yb�kB�t"�L�!��PU��ׄP�CP�m���4N���eH����D��Z�4�������>����%��n����<~ T���2�p*%kĭ�ГѪ3P���%�\��W9*_�}�U��{'cA"�w�����9k�v�����@��u�ڡ"�;�G����Gy���t���<�<��iۖ��@ФqK��fqx�"��b�a�>8	!�D�@
��"�P���I�|;���'��hK�QcR*��r�����SgNq��)VWV4��8��6��j���`��8��)SׁS�N��K/s��T�g܎��F}�9�"?�ϊ;}V,0j�$3�v:�A>� �l-��W�*��V���He-��r&vjN�6C�M�4̈́�'O������E�f�~zp���� =�1 I�'V%T�␮W�zLU=t��h�����!��".����x�P��>��g�(�7%�?6��4��҉�Z�Y<��Ef��i��0u�Kv��w��P��7����nv`�S�#�6�-=,5��Y������f��
YmEi���1v���eN�9é�'YZ\"Z��$��f�Q�
2�s��K�삞&�q������`�c�"8穫@Uj�`��l��)3�����S�O��ݷ����g��Z�`�7���R�b&�7��؏E;w���v�ӧOs��)5ӛ��Zt��~��D� z�
_UTe~ˌ1�)mwW_�9�|e����=y���0�W��|v�QH#Y�h3��u�����q��Y�>�<KK���G2���ze���9kΪ��*̄��M;Ǟ�#3c����|o�g�w�F��W��VN�(��g���"a?���dM8�Y��B s��M�ԷL��6b�rI��(�f��^^��?�=�fB}V�3'��9�	J���2go�sK��,��䐒�c���ç�=,@�q!��3�2.8���y��9���pX��3Ŋ���~�(�������},��Zex�q�l���?ɶ��!C�r&�h��Z1_��Z�����#"Z��e!��ٳg9q��!�i@Q���"�	���<�QW^��N'�X_���IN���W�wf��X����D�R��e�.#x4�4Y���F7�2����+�I�fj��l9'� �VtJ���%�r�K�AA5����~�K�K�u՗J��1�\���&Z�*a�6I-;�?4�f�;Q�V�:��g��A?	�S��km{��S�S�U�F�[�|�:\ʐ�
�`U����h��<6�I�EB�x�99�D��{��ԏ�=��a&��3�[�rh����5mK����Ps�B���ke�b����I�O,����j�����*�_8���*aP+w,��4�IAi��6�P��*Gۣm����.�4ThI!*N���g=��l�gi�L;������eV������F�T��d�FS��7�\	9TU����'O���:���� �`���Q*e�jA�9��N�s��uĂ��
��}�!�����q�@��a���
�KK�C�T�+|E��@��Jͩ�V_{ߺ3�z�w��>ۊsC��4X�@�Z��k�`0Т��3F��1�����I�	*"�������ʽhʜU�.�A8Д
)�u�Wӟ�v��N��q<�0���M9e
Z)�D-j�J0\?2��+Ѡl4A��+�_���e�N�� ����*�Jz��ʜD�"��ӣ����t�?�3
�������Rv��e�)���.#��v�1j_��5�<����༲̄Y1�eZ!Z��@F��s*�Wq��i�>�<ϝ}�(y$N5��^�����`��^��'s��a�T�A��Z�Hs$uM�OI�x�l�6N���������� GƋ�9�"�q|��kA�yf�PP�8@���Nk_A.�eF���)�Ws���ȏ�8�������%h�������7])��z��0���1mź9kc �@�r�9�	������fE�i�j�(<���s{���v���S�Q��~���J�ٰ�g5�	B��e-B{ nfn��r������SĠ�d�6�#8G������RMk�$X!3ayy����f�Q�=Z�"�o��dJ��e���pJ0�B]������I��Vg����WJ�j�*ЙR">��6�@6�A��r�j�Y�}��}AUq�e�8LPʺ��~�C����ams�*��F�K�:������q,Ⱥ6�|Щ�Sq�R~\pƊ�߷���+̯����T��7(�����S��3I.[��3L��B}B��O{]:��֥U�b ��
q7�C�L�ޅ�g!�}���9ЍU���ٖ>�t����?	�Vw;+1������ �F�8����ΞHͼ���e>d�慐�)E�?
\	�R��D�Q��^����BׯzB���[c��ᐕ���@02]��7Ηy��aV�9uv6Y�K$[�p"u	DX\\dqqՇ�T���z��������8x?n��y,��ڗwb2N���"���$淜�����[RD+>C���Ó�V%�۷�phP_�� (ͦU�.�% b%�{�>�̼>	о��g��w��}<�%�礜
�L�r�d��Tw��
*)G�3��[������JY���ӥ?.8���>r�y_̏�8Q6��i�uCe���%�R�vjPE+�HS�v^y�H����7l�9t X��1p�$4�:vj��s:��ґt< ؑ3d-�~Ф��0��m�c����;%���HtQ)H��w�I�CR6�Ӓ�S$Yy�Lo��������FL�.��(��DZ-\�!�Zhw")G]�l�ֶ%�R��PK�i��B�
Q.������gQa�Ⱥ��6>�Y躈GUUx�13��gA%��Rd�'h7r�f�*����ư����,���n�g��7edR�j�Kp�:u�����,�`�{ �QgGU��T�š�
��v�	:���uJ�%f�Z�W�̢}R���L���G�c��?Oz�S6Ä�ٳ���I�]'�愽�8f���k����~����������q�����<�?ҍ�A�H�K��+���B��?gM�E�D{��~ڋ*�T�t�հ5
�V��ߗ��3YE�ٶZ�b��U�q�i�F��:z�5��\��J��S�N�
�*H���]��s���A E<�kf��i[-qv_+*�g����I�cqX���`%鄔2��.K)Zq�������������B&�1f��(L5��\QJ��kbx�0|��4�����X�D���~Z9�Y�YX[]caa�:}�$�����2�hvH֌3�M1�0}�@�6�>�0�CAz���I�W�����O�)h�#����;�ؒ����1�3�;���0�#����C�{�����c�SR}N�($���'#A��z�9�Wٹ�jO2�c���=A� I�
��R4��}�8o��]:@Z�h�e�41���iZ� Q��aA��
Aˈ�4$�8�}ro0������,�w�2�ǧ$��г����Ҳ�f�T��K~�Q;ʎe(�d�/tn�wTD����Q�@���"m�O; G~p8uzy������k)�Z��j��ڳ��Ġ��P���9c��G�+8�QͮC?ro�*\*�=����?l�w���,SӍ�6�����9�����'�_��2�'��a�{��P�R�a���ٗ<���4?3���\"Z�-�4�/;s�Xdi�~��$h��,9���4�9
S�T4^�Y�_�vB��!�T������M�K̔�4��
c�g��K*����2�������!y�Z�i��,���'�bg,�JP��5�~�m��!%�%m�Q�I�l�DrIK�=أ{��w��m���<x�u4';jǙd%���Ҡ,j��3>��A��3���a^����`��tW��Mu��?e�6\9k5qb��D�:ec2%��u	$z� j&ҹ?�γhl�\C�-fH�1���U�Q�]��㠅곔@f��B�lm�i�ǚ��Drz�|�FA��ggao[M�`�5��qz�.�]f�rS�w��o��
!R��}���m��z`��{>2��O�������V,��>�u>�IAF���A�Iھ-	��4+s �����O�8��L!|�}�d�R��D?x��$�85pD,�D��W�&�j]�	<ɘyX?�i�E�"bm�J�j�t�#FM��>A�Z��el^��emԲ�'w�6�SK���")j��}���F�hS������e=�:�R����ǖ��.��H�z)[�)=OYs���
���2�0(Z��P�S�"2����F2�i%�Lg��=_���Ѿ9��M�8l���^�LBߡYd�2��Mq�Zz�2_��T�ŗ5������ﭞ�#��Yt>����\��~9�* X���y�Q��2�Zf�)-�η�=�~6g�zǆ'`�~��]�x�J8��n�7���j�H#]��5m�9b�&��ZRmʜUz�!�Ns����4 :���k-��R�W��I�Б�~�Uc"g�L�dZ��m��IF����@��A�R�
����T�#e�W|sT��F�<ٌ�#��C�2�Շ��dk~�5Ju��c"�iE"	IB�uL&�N{y��e1��3���2[]ߤ��}6c&���/4)~�J����+d�L�S�Yl�?�S{��#��H4�IÀfsj�П�ܵ�������a2�h�p�@4��}p��<�n��ݤ�ě�che����>�4�VџH� ����-g*6�Wz� O�R�&+�䨫���"��,����K�,/����E�XZ\bqq���e��[Xd8���a^͉�'�嬦��M�fK��$3��ZZ-��W*���0�|�y��R/��TA��h�z (��f�맮�H���d\�䬜�hH�1	���RG�u% �{�>�9%:P��a(�j#�-N&-��#���t�L�n���x#=�ҘH4�y�s��u}�N�R{�$i�R��\"�bb&==��pL�2�U��D�!~�h�VB���.��i�,�}��#��B��^m��+}�`Zc̙$�h�n$'R����><����9k6 @�F��pq���e����'�7��8���)N�:���g�ƩS�:��?O�dcc�յ��p>�R��"1��C��Hf
�� �����L�#��:53�҆�i>H�Z�f�H��n)�Ź ��:̨H23b�]ך9.��l�@.̪��G�Dl:M�/�sOu-��Q��K��#w�F��-�������#���h'bL��r	�������	<�r̴m�x4f<3�hK����;)���l�U34��{(<�#��QFF�0g�vJ�YT ��O)BJ�ց�����x<�k���P@Ċ��R����/H�[����ְ����O��q*��q�p}��:.�睷��>�W��%���/�~���/>������|~������|�����/��˗/s���YX\$8G��d˫ߦ�?*�i�
Y	�����p�:Rۑ��R��ɹoCM�T+k#)6��1/�o��Em���}�R��'���r��]vF�����I���-5)&q�4�&"��i���<�h�^7�#�hsd�u���rм��@[�5M���6��ݣi[5��\v���V��Lѩ��m[�v��w�wo߶ ���4Kb�ҜE�H�Oqj�k�޵���,����+H��Eö$\R��C�+��S�o	�(pws��F�Y���d5v�p�MȨ���A�U�w��O�}�^`��,��������]���y�O �#T">|����u`m}��.����λ�������o�?�|�7�|���~��޴��[���ۼ��ۼ��;���ۼ�λ��g����o��+�p��i�C�h�|���Y,��h����,@E�@�dڰj�ZIF�xΑd�a��Ę�ZK�=�(ê�=z�[D=���;��tQ�ɅHZ`�U��]/�ɪ��Վ��]��A���M����n�fo{�6i�RB�ƮT�]"&�����y����cL]S����QM�]ב���u�v�*�$�,�vZ	'B۩@���Mۚ�Y��rZ�D[;�)�ZԬ��NJ�Վ��=6�6���E�&�\j�(sLBg�R�H�&���%�r����{AS�~R	$*�E��J`U��?�D]jIm��VN� -��п���̙n2��{lmn���o�Aǡd��̉�5�Ct�T8��3r��N�QcAZ%0�1�1�5��|3�芦v��tv6���v���.�4{���s�xn�d�A�����U������Ν��ƿ����������孷ޘ���;���{o���������g?����g|�����/?���9��~��_���%���_��_�/��+++HpĔp^C*r�5��2ǧ3���-$�Hđ�l�rr��%�DК�1F$G�<�D�����l��~�}������D�:R�H]đ�9B��b�PA���J@F9Z���� �k��?PG!���VL��eww�[�o3���u����.��n�Q��Z����Ѭkk��MP!��!�����XjR��T'�`z���x��Ύ�U�S̤�z���#�iCY>�S3�֜�#{{{����s֟�]5�XN_���Uc� �ì!9+'��$�g{p�֙�"ԇR�!'R��]J�x�Z�Z�sd/�icd��=�mn���C��.<}mJz��J����#���K,9����GL�,Wy�t�Rf[��Tk���Y=j�_�J��o�yp/�gX>����p?����Ñ�3j��q�p9�8���ʥ���t�"gΜfg��QG�d:���u(3M�0ޛ�3�a{k���=6�����g���do�xg�xw���]p�3�N��+�9w��'("	�BJ��|{
CK$mJK>�P������N%:�αv�$ykǉء�vB[�+��r~�NQu~bS(h��"��jt��i�IM��Ё�_��3����¶Y��"�������P�)`��E�ܽ˗����6I���*�{��l��yf�4µk�]�B�2sB���-l��Y�Rl[&M$�	1wx_r������d�KT!�4�7nr��-nݺ��:#[��<h�"p�ox6�:e�`�Q��������s�6�i����!+N�At	5�˴1�ִ+���4r9�7[�I���r�9"���ض�mK��/��#���2j�֯i�XL����-�ܻ������^�N9�=���{�︠+i�s���Q�� ���ڮ��Rrx�+e�o�Oq� 3�}�*r��&-��H��Ҟ��<n.��=��Q�ٛ���!Kv�׾f����8q��_�̙S���3i���I$�3-�g��HDR���?'�,\�����U^8��ϟ���:��E��G�>�~j#�C���Ab�|�&�X�C��;)Q�l&Ԯk�R�tf��J�=��%1Ϟx��}$k�Cl[ڮ!����j͘�S3�]L��{�9~�9�W9YG��63((���w�v�~�:�o�akk�r9[���}O¶��]���Q�1�1w�7AǾ7��[@E��HuJ�fN�^{ܴt͘6f j�wV���i#V�V�����7np��-vv�տ����^���b�MGg�3�����������[ܾ}���]- ��;R|�Np�tNqt��c��tڑDr����[��=t���:܇��C�@n:�fBӵеD'Hꬭ�I�����1j���m�߸���7��z�(x3y۟�@O�l!ϱ�yВQ�V�iM��ttQ�P�9Y��V){�0O�ɜI1�6m���9N5w�v�\��BU�he����_���)�5�#g���O�s�����Ἒ�D�	�Ɠ��^�h��5���6�^(��掶i�[�D)K��N�����Y?�N(�!h�T��O��ã��+Lc���S\���R���4MC3i�����	�8�Im�QKR��i�4��8V�0��'gmgիc��f=˛<|���{�?s�6�Wo�N�f>��d<bss��7nr��v��h���i/K<b�X-�BȤ�е��d��ւ�}PG��rg>J�"�$-\�#�IK�N؟�I]�$gmTM���+�$j�����^����w��Ыc�!���Á��2K�x�Fl޽���׹w�m;�}!8��13�(�L�2��uKil]�1M1y�i*	�,�>��(���#M��Gt���A)fi��(K��]�жRLܸ}�+W���w߲��Oj�olէ��N�.�S���H}��uɚңiR���t�}Mx8{�}��.g�vBӴ4͘n���	����?d�G�<9y����a���� O]Y]]��:��kg�^'|�b]ko��K��,,������2K�K,-,�������`�T*���Dwt�!����"K���* ��� ֧̿5 �~,=�i��x8j��fǩ�11nTx�j�z���˱�]&\�Ŏ8�?ڣiR��� A[vy�'hE�~�z�B�t����!_��x�J�$4]���_|���v���}��=�,�¡ͯgW���.mj���Dy ��n^����p��Eu��C��HIH���kcj��
G���5�\��j���>W������­[�����Xk<������L�A#�d­۷��/��o��ܢ
�]�iF#�9��d}N��ڢy��y��>��,�S�"�ܴ��S�x��4�"9����h�P3�j�P�C��t-׿��W_~�͛7��W�!���������t�x�7�#�B.�m�r۶ ڠ�gd[����4�$S���J�4��uĬU�\r�T��5+�?E�{���ɿ�Qd�����
��_?x)�A= �ܶ4�E�J��U�P��2dyy��e�זYZ^�ߗWX^^fźG,.�BE7m^�5�����ì��H��t�m(��E�j���&iU�IZI$e5Y殳�֬f�9E&Y�&m�U��F%U,�nj�>0�@j%�эƌ&#F�1�IC�i4-��Cs�JI��p9�f�j�)YthR#�}��cC<�9M�p��	�ML&-׮^����p��u�I	��Z�bk�(�&Fr�%��fD�ut��i.�,Z�"�>a�4��#m�Ķ��c%v�F�O�(��-�^�%�G�h�1��͛����Ϲr�67��܎�&0G5�!8�z-�4	>'M�������믿��͛�'c��BGk~okz\"�U��r&M&Ħa<�躆.�V����SF�e���,_?"��.Ҷ�q�>�IG�K����d+��>q}4�ur1%n߼ε��q��Uvwv���'O�6�>`�d�<goo&c�9w�1ѦH�4��	m;!N&�Y�H��v�D)Cn�u�R�)%���t�qK�6�SG�ZR��
Ԓ�kӿ�4�W���R�J~,xn�=��:=$��C�����"8�O� J¹D��Օ��O����s��iN�<��3�8���Omp���l�����S���3����e:���ӄq /N=�Ԭ6{�y���㸠�Q������],W��HƇ��$R��4��n���ӂ�d�/цsS�Ӷ������}F�ml5�<�h���sVY��{B��OO�!b�k$#���^�q��W�q��5�G{d3A&�3F�DDovCo&B�����m�Դ����v��
��z
��P3��c2n�L&Z�M"����iԤ�ꪆ�Fh��kW���ǟp��5v�w��(�c�}s��?�g�8y?~��H�64.��`��x�۷���W_�ݷ߱uoK��|�wNn���{�"BL�N��m�bG3iI1�5Mi;�Ԏ�!wD�����ZU�Z��1jF���y�~~�pqY�.���U�zi��k�f·�]��k׸q�mۨO�i/��i�AH��=G���5]FR��V�6���hZ-���,ϲ�3�N��f=��D�%�&�u�ZR$&GvϜM�T��5	�7��3�YXf�@�c�<>�����P�)=��AJm۲���h�XC�D��p��;���*��K,,,0.�0X���������:,��X���ƩsgX_�@B���rN�Q�)B9@�a�Mտ.����bf��fT�.����@D��5G�i"M�cC��MC;��c��}�{{���2�1��@Z� !;�^�ܑ:��*y������VP���:�$��F|��7����嫯��7�G����Mc��,�.)�ăK���)���0n�I�d4a2��퍈�	�i���8ni�M��tc�vB۶�6"K�(���s̚��<�itn*׮\峿|�g�~ƽ{�t1R�I�Y3��K�9|%Tփ3Z4�wM������'���o�-W�x��]l5�7��s���M�zr�413��M�17L�	�d�x�0�ߓɈf�ҵ���A�{�2��}��^��ji�cB��چ�ǟ��g���k�ܾ3����G]���>�]EQK�h�ژ"1Fe�Q�]����4�M�d2f<V�v;�Nt��ɘ�m�]KgJ���&L�/���[Y������'~G�Sb�L�Tڵ-��}n޺Eی|p8*�A���
5!���W���$�*�	�P����a5d8�j��6�������$k���jq����O��ۥ��1�O��E�CI����2�~R@֜:��Ӷ��a�v4�����M&�NF�O&��c���ڧ1�T:M!�Z�=F������&�����������Nn޼ŧ�~�g�}��o�[[.Q�p�x40%f53>d�8� �%�c�m4�e2�0n�����ј�dB״��Ȥm�M����-,��]T`��Wx�����6w�n򗿨_Qͣ�6Y��B����!�![Aw��\4qD}b�o���/���O>��۴M�H3N��suq����g�&����h�	ݤ��tj>�4�mҨi{<��MZƱ#5Q�P8x�3�@�9�xRj�q�6_}�5��n޼��޾Z&�����@�wywG�t���挺p��F;3�:c����vt݄n�0)k�vZd�А��� (h�����0X��aP<��jx�w��0���S26}�G�Y������o�1n�,��*G��a��@ʑ��0�ڦ�m�F��MZ���U�������p������7o���;Ķ#e3_�|�)0.�4��A���}l�Ц�Go�2s��c���
fr5O�h�D h��3M�tm��؛L؟L�oƣ=�{c&��1;��5//[%�h�(���h\��n���HI�Q2Z����=���k>���|��Wt�}�*�CU���ZP�M�Lz���&k��.u���h<f<1nF�f<a�D��h'���B��Y�2��!P�/'0�kvF�|��7|�ч\�r���]�wT��[�~/*[���(��3��ݻw����裏���&�	++˄�%�45�@<%�6�����4�%��I�m��al���vB7Ѩ���Wv�����)�e)NZ\U����x���W_��O��W_~���1����X�G�c�'�ڞ�H�#u����i���iu��IL�c&��ۤt�j:�NM�m��tQ�����-���YKfZV��g3&yf�p��p�}�gp8������m[�����l������u���Aq^�^Հ�EN�<��y��L��"���HY�r�/a�Ѐ�������O���?s��M��ɘ&U��I$C4��!��E����F��A�ɍ���p��/���d�I�#e7f�L΂s֍��ϐM]Jy��f�E�k�}8G�����k�	�)����bLH����5Ϝ5=/%��)eՠR�i���k�\�µkWˌp�A��U=J�u~��.v��Z������5�D�Fb�	��[mJ�!�iE��|s*B��gF�܌}����@�t�û�Z��#�{1_"�O�YUݽ�=>��c~�����?���߲��G��l�0x��ȞO>)��+	hz���.ۚ��2����	)f��BP�q����j���m�=������c�h���+��� j/Z���{��^���8�����.��G���~����^��h4�smN���^)�jt\�=a�1��buu���z�W^yU=����B�w�dfʙ�A�X����������X��#&AD�i��p�y�V��	�Ш�{ތ�AG8��j6����������7Z�4#�ϣ�I���������ß\Q\4k���)'v�w�z�
�~�1��#���*������iЄX�h����Bz�f�����{5Ϧ��ވ+W���O?���?���[��G�	�O�L����Z��H��i!VKA�X	F��9���$!�8�-�|��f5Q���	�$�W� ��|��	N..�)[�n�����Ģ2�?��a�$6�Z0B52��OJ�[7o��g��o��{��џ�u�:d-�(^��Bt3Z�-'4��)�tN���-��d�������h% ��Ȣ︼g��h~��|�~�!~�!׮^ekgG��C�F��>ǃ�2�rLŪ���;F�7o��Ï>��ۿ��?����o�4BM�Z�U1\�i��ϥ8�A6��fb��hF�L��� j�!1�Py��v��˯���~ǟ?�3W�]eo�.v��b�)�ǵٚ�Z�8=~�c�^uN}�Y�gU�ԟeO���%)�e�$t.kxa�1[�������Z��h���d%.T��X[+��ڞ-34�_���ԄPh�<t}����ӆC�OA�����dj�i�	W�^����o����ܼ}�I;��QkˢR�,�� ��t��V5	��������_�������O���f�v�h����Aa��u��B&�����m��5�_�/h������!�I�9kQ�n{��-]����ə�&Zcv
�̶��*6��u���x����E��ϱ]U~/,W���<dxQeA�WY�F,���{$[;{\��k~��_�_��O?��.'�aE�uZ������������iD&�H0�mu�4
Zv��
�x��޽���G���?��>����_mv��
.T���~�ǁ�� �V2�k�=��ܻw�O?���ݿ�/��������w�P�b�D}�{=�@����� 6?����tn3�nl��e��b0p��->������>�Xf��
U��s�ܲ���g��G�σ��w��y�}I�Y����)g]/D�w�J�fC���U�2: ���1�Bi��� ���j1�VT+l����	?ٚk��I��*�th�h�O������x��9,9���д�6cfww��h�s�`��q�h5�HY�1YS����|`eu���UNl�`ay��/t�� >�C_Ӕ�,�6c
)�>�h���Zs��n ��;�eeH�4�FVB%�|C�f�/H.f���tS�����k�d-����J�	�s�|\Z�S�5`���,PY:O1�gc�nN7QM�\�':�L�����{��$]P[]�m������[���Nq
+�E�;���B���P �>��L2s���ޓ�e�����Y�}�}��}�=[�E��n�
辥�kg9cm/��,�������n��VSrd8�0*z�e�nf]|`��P����׌��3O��uގ��
�6��d*Å��XS�s}E�܋����:R��c���6�L�ߟ�R\f�^��<B^��u�����X{�"�`<Y��Y�r���!,?8����#��
p� ��2{J-�XhN���ӻT���q��m�(Og@��ys���B��'+V8f)��Z�i9V����Q�QzL�F1/'�)�~��&�n��8����{;��Ǻ<��*�ie��艃	N��)i���Ӑ6��2��%]Pp�bֶ�I�&5�NK���<���䋩H��r��6W3D�����w�ڼeT�W��<n<�bolW8}q�$�߼�SH�817��̋�"���M+'�\B��ۖ单���,%z�l��E�D��ku���������|���Ǚ���އ3t*U����@	D3�c���|���N'�?Y+z�J���������!��q���i�HM�Z�QZ*�9m8������G��F�ʋ\*s��^f$�=��h�ZI:h�e^�Ys2�],�Y.r��j��cbSo����"^ק��8b�>��!ڸ��{%)�&�C��r`2�a�ۛ6�gz���ɧC����cfݥ.�x������N�y���.��CX�Q袦9H(��2�x8�=�c��c4��9�Q*�[� ���D��3��;�k"G1լ�J@�����0��Eҭf���:�=]�A����}��kE+��u@�k�zZ�+(��d�tk.�L65������W��s����y�e2�M�T���GߎIG�Ɩ2+��j?�1�l͟�7��փ�AjD7����9p��JH:V#��<pw����7����	��i�f{}��R�q�A1�w� D��Tr���Mv/�t	����G��>�ߞmX�ŤS��6_�۫ݳ}zO�c����#���w����i���=:'��u�M;��Ty�5�6p$�X9�p7&чc��Hr���I�߇�o���Mz�td\&Y?_bɆ�	����nXKw�f^�&�G��I�aB���;�LJf4����������_h�El=%s�84c��X(4ڵ��Q���Ⱦ]����[�Q\m�b��k��C����(|������7��
b���>]9�^,��Y��O_��<d��l����sL�}������ŽM��{^�yW���x�=Y`�n���O�?L�N�����|OȺ&�/��i:�0���ϝ���+	�8�q��R��p��q����KTx��V��M
7���ݰ��[04����⵴�b2�U����,�1�cީt��z�x�Ƣ�~C�r���튂��*Ȩ���gDE,�d���nÍ��T}��Ϥ�.e����s��jx���s��n�Wfvޞ�����=@s�77K�p�������ZD6
L�4���GWv&��h*U���M��=�5^<�	�"��17��1��	�3������=>i�=���=��{���y�D���%���(����������ƶ�c�gO��Ա@V
���L#0��)������ˤ�[���ZH�,�;��\���-��},�_{��39�gX���0���p�Jotd���f�i4�g����7"�߶;�ҐJrpM�BQ_��srr�2�8��PWq�G�%Y漃�J?�ɤu���O�A&f{��q/>m�D�훁x��,��xc�r}�n}=m}:k�����e��|y��P�*�g�F�m?x��~���V��M�W�$n����y��m���̒bŎ}ű1�ټE0>'�Wp%&���`���Ci�m2�i�5��E�S��k���a����Z�{�4�i�(3�c��'����
��	�l1;o_]Cè�S��X�)P��5#}����O��="�Or��7	y�}����7�:_H��v�S"���g�f��l�����)2��֣�A�2߀��Z�Ɩ���M4���rM���ʪ��	�����'�̀GV�S���Q�w��+6)_�|;r���l��<7��օo�2��"���F��XZ�0MGɐ7����W�(.x���
�76��A�gLlb��,=��,��;s����l3j�3z��w��]��� �l߽p w���>�;Q���.�{�Z��7����j�G�|����_׬��J�5�'.�\]]=��.�oZ���ww��'�c���I֜,�@�A~��t��i��x�|}�ֻ�M�'���a�b���bO�������M�ӡ-�,�z`F��FId*ʓ������������Uᓳ���Ɓ�r�R{��C��� �!qy.��eJ��G@A	�Я�S��i�����#����x�榆з d�d���k��q0s�N/�!�.(f��;z��uF��:o��Uf��!)�nkX�-�t9E�o��l��@F.�e_�SK��ǩrN�-���A��- �n笺Ө�5�*{�p�	w������Yʩ*�OR����M6�®�{i�1��\�j�屶��:�p<st�����6�q���Pnim��o��sO jl��s��z��˱A1[��ʈƽpg
dz'��9o���
l����m�zH n�-�%�ޜ�&]|��S=P}�����ID���:�`t�l$ZXz����l�3�y�v2N'MA[�2J ��������=�ḩ��H��(<���-mnڸ�%�E����M��#^[z4Fz�S=c�и{W��Ɋ6�܄��擓�w��y�$	x\}B_}Şv��K�1�x��:��r/�:�{����r�!��6p��Y�ͭ�pQ�����m��ڽ�􋵦��SC��o`IN=6�xF�V�����pځ�O���7,�����i������]ӧ���w��u��΅�	tV���A��"���?y��G�S�3��O��KVc�,�{�4�]�#[�x	��ќ��UX�ֈYDG���������m�+���/���8I����[/p�4^��v�/�o����'һ��3[��g����2���ޡ� �ׯ������*���W%�\�g���,�T�Ja�s���غ	}}�|�����[��.YД�֑H���`�����}����/�'x���4�:����Ћ��,�h����EQ��G��a�Oi�߬�|������J%9e�	��f!���uw�e�˝eU�yNKi��^�\W���b������~6�ep��5c��Q���z?xN1��>���,/B�^��7|%ir2|�V~A������Ȟd���ꎖ��k���\3+�ġ��;�ys7���S���ހg����73�ko�u�1!�'[�m����u�NX�yNI��P��s��kr��:*�VO^���H���V�w9�m|\U[�fn��cO�3�pt�ޛ��u��Qsޣ3,���gl�������>�}�|��1tB�������Q�T	q�m6��.�s����uu>�%rS\���[����i��>�>0�W�Z)��?ѕ��HS,�F�%������c�s��b
��/:�O�R\>��FOT+)���^Ip?�K���� ��<�/��	wS[��}z=�3���#�o�|��=��H.�N3	�G)h¸QCG�hem���9��H|��~���M7ñ�{�cigPS�}v�����7z��E3�B�{����I�p�s���u�O���x���麗�l�~�����9g�m��:��?�A�d�����ra��* �Zfq�+�TL0����74�^�p)V*�~�]|o����bZX:9ů��{x���3���p��9I�3/���׊~z�L1�ٺj��ݭU*���]����������z���FF����8��o����I���*?�/Z~���x�Kd�l��27�e�������9�Ye�/���d�r�����
��W��'���^�hl&?b��&iJo(�Y�p��_	��ש�&	K_P���}�!=�qo�/�_&	�q����F�,�{rp��L�m�� ��� �s �`�W@r2�Ȼ1���+��"(0���)�3�p%�I>ǨtnN�7yr��<��I���X������j���ݑ��g�_ט&ڈk���v6�k��������s}c�'��N�$�3�$�n���1��5������4nn�g���))'&Ӛm��`��ZQ���e7�r��9}��k�N��d�gi&�Z�] ׻.aq�bU0��}6^��puF�a����N�a�VP����n�)�_b�#�^�6�B�<�)�[��C��-"��ۄ�93�dV�aig�����c�0M���v���ۦ~d<w6��ϱW�`M��2i��2lz���ʩ��'�\6�0k̹�ɽ�N�e�K��D�!�P��扙��ؿ-D�M'�
�mp,��T��WPֱ*%�悬o�@ɵ��Hoƍ� V��*�f�(� ��f�6n�tr����{��~A�YyaM=�8��^��L�DI�x@f�!k���ƌ���c ��]���(T�I��?|`��"c'"b@�7�����֬��86!*FY�:_��Q���I���\˟���#Ǐ
D�s������ǔx�[���_�O�&��Z��$0��5�Z��I�`�|���\&��tRbV����	W�л7�4$P��/�(&O�����Uu�=�J�D�K"l���r���r�~�g
�������
�-��]cD�A���Jf7����8"
�傋���{1��cK��㼝���u�(8��P�>+�C����5�Z�mA�Ү����U�ɓ:hG[���x��`O�� ��W������&�^c�AL��Tl��&	RI���-�5��5o�9���ސC�������>���GqwP:��P��m�����^� 3N��x)�X|��#�W�,��ӿP�~m8���✟�.�%�$�/�R�\Ip�^m��`���Wx�v0�{�.��.�tH�3\U���*��J[�7������b1��ky�8d�*�#�}��~������
&�X5p�$6f��q�.R�aJ�u1��'�Bެk/����%bmt�I�Z�K���=&����P��g��tTa�����|��H�2m7O�U\��AN��Y�݆nn�b	�JJ�G	~�J��7�����E8M�(a7,Wr2HC���~��n�~�]�������,�*���u��l��]L���J�����H��92���-���m�<ǽ��2@i��R?7"^>�l���V�$:Ֆ}iS�i��Br�bꄨ���u��Z9�՝N�}��*r[ʌ�#	ZO�&�4�]��I�䰥e� ���8�r�'9���+�JMr���<^i?Vв=�E�P�M�!��N�7N��iלj�����)Rn�/sy�l�ZM*�.���A}�^�9�j|j��W�FҠa�e�<i���:���f�q	�ƥ�1Ӄwcva�%>�[��CQ>��;�Q�.g"xM��R��j�S]�/`<�H�܀�b����LCʠ���J̹]��W���|�؞�B��>N��h��F�9�)]����~c�t�&�A�q����\�W[.��vL��qR�d���NM���s<=�Ɍ��O�r~�N\�Kd�7u�"m�t2L�-�>r}��@c�)\|/���6k�:�#v�\{���_��^D�1!� �[qV��,�K��A���`���7'��e�ӧ�
��_1˫'��@U�E��V���� m�YT�ӥ�K&��=���{�S�r$�<�|�]��t��]�*d�w�X�B��N����_�hH����^�O�%e}k*�,��`��t�h1ZO�pJ���c�����ᯙݩ�V]���rT��1',��i��v��[am�b������Ʋ�К��� o�)��½y���!��cZ���e�}rK̋c��&<��*�~�������Sk�S�������?(Q�os1��sC�1����DH���d�����d��y�0��u����/ts^$SSŮ]�+�}Waxu�x�>?��( �3�␋ϐ�]Dm�_��2 �Ё/����k�l�qY}�0�j3�?W'�#Wx��/'Uj�7d>>}<�Z��t#�X��x���+0ޘ-�?p�K�bL��.�Fg�f�"�3��w%Ī�U#�{	� �k�>��9?JhT��o��d�4�/LV6a����_}s���B����ɯ�Ma&/,~:�r&�#���|��?K���5�5?��3u�.�䢲�D�;��1�˟�ʙ�^6�Swe���*�3"�Ɠ�C6�$,\�����w	�S�����?���P�wr۩���_6���(Eg�R����q?���Q���g���Hr������FF��Sp�?}F�v��Tx�@�PZ��zVt����	��`��o��7M��Y��}�/ۢ�<	��*M�8i]��y�Uzة�v���p���E�)>���p���oRVs�L��,U@wᗝ��R+��0�ԋ�ڞ����B ��A��W���ލ�1w����g�	�0�udo�˾�^�&m��@w�*��dF�o���s�	{�t���3I�Y�X����$�������ʃ���X���vwTA>�z7&j�B���Mr�M�>d�`��^��� ̎�fS���	q/{�%C��*�u�%��<;�YY�@]��L�m���q��
�u)�B��a�rR�Y�&��o����������ݝb���h0;����8:��b����� <�+**n��M�3�?���=G��4�#2I"�?)�:%C�@Xx�U�V|�����=߆{M�Bq��'�(o�o�r��� "�L��F�DA.;7�tR�E,ɡ��^`����E�^����}�=��a��`� p]Xݓ;����kpAg.�����+�"�r�șS^a�� �nI���˙��(��=�#yE>��T���m@i2T4�|ѷ+v�%����O�\�Ȃ^���o1A!6�p�͍iܸB��E	ښ�b�������0$YT?_l��G��8��J 2��fԉy�|��h����B��'�1�1��y�_!�U���[OU����wj�m[ѓ=;���w���NnY-j���o�D��-.r�|�y0=|�p�Is�Ru?`�9/��r�pJ��t1 lwa��.�Z��TAq�V&���/����;`�W8�l��UT��b,�2��&���|�z�?���_No{�����O��зk��j�V�:��{�#?K?��E<���s��p����8��"���(v:>yN�C῁���t�1������m?��]5��ۧY]����k_�KN .�2UB3�gP� ����t�q�*�����z���ѡ�ü�_��c��A���4:���	�\4�ަ�4�(gE����	��+V�C���`�_�R����i��x��["3=2�Y�����ҝZuZᲔ����3Tm��q�Dk�-�p+�ƺ ��w�����Y�ɭ� >�AB���#���1�J@���i����G��}����]�q���f~����{CC�4�J04Y.jy�n}���SD��*�y����Ug�A �dq�P�4��IQ|� ���ܢ$&�I#�Sٻ�9�*f_�����p6�;��[EW?_���ۤ�����;zL�"���vs$%�$z0=�s����2��YY=$|*�I�e+�?Hӆ��8myI`dg���'=�W����K1���n����j^���p��|9���HS܆�az���m��G,���T��+��?���~�ׄJ8�>�I�ē�����C6�_�A8��F]w%�]�9�*��Ŵ�k���q���C3������s�̜�]]�{���4��q7=c}�����*|���g��U��$�>����9f&|�~k��^.<�/\�y�o�]J�[�^� ���a�_�f�o�;|�JNF�W��!��Q�����	:Y/`D�{�񶣹�|���$��{wP邥/8a�i��̐�*/O�%�텊���x|*u-_aT�S�W6��,jN��������Awv_��*���P�V-j�-/��T�?���d�)k�����;
˔�@l)$�_ZY)�#q�7���Ҥݗ;�Q.>n�i'�Y���Q��H�8gae�0ϞO��5�.3$���?% ���)F;�a
�c�/��x��E�W%���S�-z3�Ǯ����n����.p�n��I!��"�#�_�gXU�J6�G�t�W�?�*�1��3�@cE�8e�U:���"�΄W)~;Be���e�@��K�-ԣ����,��!RU�~�P���W���-�/}��?r14��d�ad3� R�����/���1*U ��Q�*ݮ�h�au.�J���cr�r
���ݫ7�,P����M���_�'m�}��e��M��!Jغ)��,ہS��E��wU/����o�on/L���xg��C�w����X�˟A7����5]�T`N�`׭ ϛ��%��L�y8"Ϟ����h�}L��y�
Vt�O���b64}G+d���C�S�2BM����"m&�+R A"3��$MU*��)�ȶK�����kHa��*Ȑ�GUm�
 P��Ň��Y0���)��J�p���u �nX@v�1� m-�������X����`�����O�)N�����[;'���;;�<<�VI�;;��lӺ�Eodi�g�ܷB"uݾ�D�k~�,���gws�۴ň�E�-���K���J��w#0B\�ߋ�
��:dq�d0N��X���h�
z:[zn�ʌe�ج���T��Z������K�E�>_���9�*Q�SR ��[��|N�+�m>���o�}�]E�L���b,�$�L�-���$/D��AX�Ԁ<6�儡*g��%��8��Kh��)�&�s�̑0����)�
Y}g����/_���������,��z�˘�U�/5g[�����,��	k7ԅ+�`�FIg�͂B�r}.�>::�ElٸȚhM�c9Kv�|���|� ���8
����nL���N%Î`!�u���Yy��U:�1�]11�Z���fyA;r-ds;�`�K�
�c���-W����$��נw'{B�*n5�Ɗ`��f�`*�❧-��
Q~adF�Pl?G���)��Ye�1�Ă��C��:�4����(>��ݾlNn������89��й0����0Ȳ����&wv����Y�Y���$�1m;awQE���FWR#e�j$1�X[	0�H8�$��o���X�ل��b��f��`���(G~�6�M�!��Kˊl���/b������X+%}S�����y���0�*2�$��f�u��G8�u��cL��3�k�-���=v�XT�n��b��Ji�h�\�Y0d�%�t"΋�tY|("G-;"���
��/ E�юB��-�!�@��X��X�����C��3�m)���"�p��G>�J����[�4���$`�b9��vє\�_��@
,�ٰ�D@´ۭ���H֒e���.�����xT�I�}3�+ev~���<��\v��0�'�>���Õ1o�� �ʩ����-��6�%.�+����v��GPg��Y�[��Čr�p��s��:��U�hj�'Lʨyj`�ʢ��Q���>�bO��7����s����_#��u�%���}�c5х��s"D�X(��&"�V��~QXM�
�m?Б����8������_F���.�����.���͍6�rƴ�O��JK6�qg[��ۨ�hE1�	C�q����6eRt�Y���v��M�J�>�.��$Y��;�^�M���-MƊ�oG�J�Ję#�������A AD��g= ���ѣ�~f1k����Jx�����*T~G�pG�\�	K�ٖ�Y=\_y�9�T��Wk�Ͽ_�
��Z� �_�(Iv��?��r�-�l��TF# e�,4��s�1���䨄s����G]�p�u<W��2��	�~=��:���ȭ�Nv��)^�D]�>���9K/w��5P���o�.�Ƴ�;��ٌ;ş.)ڞ썼�E
��%y�WT��28��H<7�e�}�i�IU}y�	�fm�w�e���3�mΔ��C��.1�C����#��"%���w+9a��4��g��@�On�Z��8���;;��dzF3�M<�T"�d��X�$vc�}�n�|�gN�iӶ�oɹ�G$),�t��I�4F=B�_O�Z��:�.)��F@&��m�����7!��ˉ�J��H$	+�ɔGm�Pk#V(���r��8.m,�w�^mur{<#ー��Iu��/�'�'J98g����Y�A"|@$���s��
�t�-,,B���LM-ܭR����*���yj��:�F�޿����r<[�X��||�1�w���U\գ:����뭒�]��i����$�ׇY�h�r	�������7s�~�\�X����6������X�+'i��䨀�^���mF̰��t�_wic���)�Z8�[e4j#>��a&�GS���-ncqxxr�L�.p���Ռd��G��\t�0��
S$`w�.�+610(�8�[��.GG#WcT6M�c�.j�~5VYkw�r�1ڃ���v�,.o,��u�8~��~~�#@:�O Eb#<8�K��Ϧ�$���jB��Zrbf��T5w��>io�]ss ��x{�57��P�i��	V
��g��d��ŷ�C�W���[['�+nV��]��c�q�l�4
�Q�D�����>�z��x�����&wB�d���ڋ��B�+D8�D��A��������/q�YX��,�[�M}(#EU�WlL0k��V������g��]no��u�Ld��Y�W�!�b�N�܁�Ty�^���mt�y��I�����sE�=�@�I��e0�򩽱���p�m�ә,l�U'ŷ�<M�MƖo\v���T��ǖ����������]��*0�juS���R5��B�$�_�OI�rx��:����`� �Q�s���Q��dI�
@��m2{��=������ <?������K�v��@�����x_&v��A�񁆥�M.��:c�=[�]�6��]�\��N��峳@A�BZTC<S��HJ_�v�-�%��\;w��À�Ҕ{[H��-��X�����E�`W.�1۫�?����t(������}��km��$�1�+s	ɘ]|ײT�P�ӲSM9�2@I��Z�c��oH��V���{*	�������"A�ס�¢�����f�nY0f2&K:]A�|�C�6vbI�	�y�m�vs+˩g?��G��
d��陡l2.��ﲜ?¢��nrxI��QG!'hR��!���� ����wg���_�y�������G$؝;DӉ���ί�*������q������A�l=~vƶ��?�z���8H��o�Ş=к���㬒A6�>�9�2A��P4�ۨ-��y�� �PV�����Β�������P�Q�W�^1>>��o�r�p(oH_
.�@�).F�cr���o��éC}o��z�r�q��T���*��͂}};���$O/��\�侐4��Ք�MLf�XC��yz���	�`�m䢊n�2�tVkl��Ee��C��~�\* 3oym|xx��CQ*5A���Ez�̸,%X���	d��S���z�����ڞG�o?����JdO�>�e��B�ƨeZ:����!��W�R��,���v)����ί���et�6�24�HzU��]j׵=����ۊ����͞�&����0�+-ӂ��#�Wf.�ns��G�I��1;��}
����l�/�F��x_�\Ș��[���%����	rl��˕rSX��M`xG̶_��L�:����:尗zZ��I6/�	L/��{��g�>�fee��>F`\�RS�6d��}�/���G�.�W&���Q8F}�W����U�PU]�F��6|���y�L|����==����ir�,�zuVm�an^�x�l��D0"j8^�a�_Pv���w�����?���!��߹2�T���1~nu��i|�Gu�Uz��.�@�gVN~��6�C����w��07��5����U��-3No�p� �lvF�w!��Am]�s0���e���C,����a�Y��NO�Oت�YCw�⑔��.�T��$�#�����c�����Y��(�FL��-��B�~��3���	�-��sA��}��f��WMC�v��X�Ҕt�Ԡ��\��`���%�BƱ���-g�W<�76�ukMv�����'���i�u������PE�p(�U,Ȑ�YＯ7�@�߽��p�(��}bVV�%�8*2�?VT$ƪ�0���M#���]��g���?��e�3�c�T]���B0��#���A�����&��o��륽��`Wd*":�(�O��F��4|;đqVWa��K!�T)���c�i�Z�k�֜h1���{�6���I��b8��ŝ��WP���e�$wi����}y�`a��G][��e7�w!3����v��w)kww8�RT��Ǐ��~ja�͑Lu:*��}����-���`�֓��6�G6���1��ɪb۫��.����!��ů�5����Q.�Me��9oI<'�L�����ͤ�o
�����⊅��lK�'<�Ay�'��F�DR��#���j���G���6|Y�˛�{g��~��~i�w�c��}�����]��鈥W����.�6b ��X<����˯^�x��ｹ�=�Q[�C�o�!_�դ�j�����>^�т��9� &��������[&��I���z?fڳ��}_�[�{/��'ޕ�fѷN�f�ih�Jw  
P ~�8x�s_8�~5(�-��5I϶���&\;Ğ��0~Xi�W���@��*1�.���L��4q֯���&��E�`�'�
N9�A
����!������?c���~�C��:*�w��L�5/���=7�/�Ӽ���U���4�^>�W8��4 ~�X�:���l�������oi����c�)a]Gpt��7��IA�=���Qv���p��ߔ�<��8����(�� +�w�`������>§����m���n��Y���#`�����]���EC�UvW��:�7l0�Q��R0�6`�����Iw;������(W��+�� ��"g�R�a_���Us_�/�~V��]�VD����D�_ �j���M����0��%�|d�<EIV�(���ba����}>uK���V�V,�f��JX��*�����?3���c�~��	�ZZIq���{�h<�#khg#`���$�&��"H��
N������aC��wA��F}cc�cT��{eQ�>�����tTTb�\L�dB����2/���<򺺺��X��i���	�;�x���R"����JAMS0�/����:qIn���]$�Otݗ3�!�0"����hkoKUa{(d��P�f� |Caى(��,MDT�`S�Դ��1�b���e|
�������c�iRxxJ3�D���{�/k$��P�7�"B�T��S=[[Hy���{�Q��~ =���۠�!sP!�Q�WH����P�$��쌓8vy��FIʦ6Sg[�H���P}ѽ��w7=�Nb�$�6�8��$��*��n��Ʃ��#.ˋ����n�v�<��M��!.ntuJ���cX9��,/g��Q�b�5��;2�1�
k��~;�1�"j�|#�䌻��1�W��s��)���j��L3�_rm�u|��Y`C@Y���H�/z�K5���|a�q�GN:4�R�&�#ftT���J�O^T��e�+H �>g�g�c����i�A��w��(��+�EVA{fv*i�EN����f��}��C�[K�LmM��s��/�\��J�S����G��!�Мz=�f.���2-M���2��nv��.�nWB��D͎D0��Ge�Y%�r{Ā��h ���e�-�6S��Y8�_�y#�GNS&�pw��Q��ח��'��].T:p�F�U��|�d����.k�s� �{O�-�����o%i��k��R�9�%���+P?��k�%V�N:^:gDc���о{7������S��_Oop��]��LB'~�Ԡ�l��\ �wC$�>�����������~r9��A��?:>jF�aU{������\�2����:�mc镀��U9���?�x�z|��-���?)��wM;�>����t=nt��`,0La7�<u	�Z!/G0����waRwAn3����`��ϔ|-Ɂ�QK,רl���zzf��S!�/���:�)��I�q_c�fB6&����x����u{n��U�n�����m�H��}n�My��;à|7N-���y���?kQ�OC��sؙ�2��*s�D���Vٚ����Ie�o���d����`����6B�R�d�|~T��pb83+X�g���rv�,�Gg��[6�ݘ=�e�����z��I��M�ݾZY�f���r� �j>�0�X1�?V�0*,���Xc�Ȫ�'^c��l��\�jjꛚ���J��Ųb����2	�(e�aF�����W\��y��(�/�2��sr���#Mz����ı3��E�6�FN�������7�m'���@�O $_��w~/#����������͍&`��j
U�|�#7��4<��1�Vz��uy. ;�����=�P��9����-��'���~�D�j�(7)KCCC�����'�<9�>�>哩jC���p/�g�+G���%.{�5�����wWۤ늋9�RIHyI�:o��ߜ>n>�&s�]�QЌ-�!��$q���f�Dy�%�߉'���,�l�-�Գ*���v�h�ߚ�����B&�%�;0"���������C��!S3w�0����f�lݫl�~5�TB�#M�iX>����6YқRX��3��;�Tu�8�tvg�}Q�
��*X���>;ٝ�]�c��d�"��>��[�b��эz�2L�;��s��$s/�j�N�/��/BGyL��G�$��֔&'��_��_[���V��"�}6�����>m�WyU�-���IX��n����
���g�����o{���<�aT�wp��t�+g{0z�+��+�H����̇�e����4eD��vQG����{C�=��S�����|;g�h�0�P$��Y���V�����:�,(�M�2��{��Zx���B���`ͦO�!���5�K��h�~z||�q,�.5.ms�[�oSc;��`�"��Ҿ�j��C��l���4B6XV�:5�X �(nc���M(a=$��H�4D�Ri���K��X���4�+������(�4ۑ�Iy�0�VWu"�&b6S�b����eag�H`��f���/߃d�t��3.�oT-L$mQj��U<8��l�S����?
x��Tb9�6��aq�;i��G'�6����&���յ�5�8a#:��&���`yV�dOjUd������8 �c�������_w_�G�g�` �g�K������s������ʌX�%�E�c��&*S5f���B��$��F�6���ľ�k].�p��Vym��f�Ǹ�éF�0eiq|����n�֓M$�xw̥2�77HZ�<�Q�\Uc����У{���$=g�27.�6������[��U�.���j��ji*�]^������NK"���c�)W2���"u��p��El�"��]94~%�V���\��,A��r��t�ߒ��e]�=v}��7h:o��Ae�*�[d��]dKM�B=/�c�d!�g�R�*+38R����wt_la},���sV�&�/����^$Ϸ��v��T!;��'��@	V��y�轧{��]��MoEMڣ��8\�L��d,�#d���O�rh5���b�P��@{� ��=�ݠ>0n�2���6c���4�Q&�^/a̸���l=s@ZJl�u��]��s�[���	�����,)���}�������@\n�ݚڛ�4Y<<�4�ԶS��d��b�YK>���m戦����*��KH �%kgM:&#Y����������_{_n!��'���ꟷ�d�o­�6&�	D��V}8�5��M�kS�`��RJqA��p��{?�.�ͳ�����Q�C�q-�����/�+D�`]�Ҍ��B#M��eIg��O�dr.�Q*�tS_���'�9�o*�H,�v�k5�M�@7|�%��8�q�h��8��<B.o���7YN��sm���Z��J�#��Ҽ�������QS�����^x�jC��v��+�����~Y�0����uD����l]�);:�N��VZ�
--�� �@9������a�쐑zC�L��,d�y�����p������寸p��+��]��Z�
]&$��ɊD�"�Z1r���1r�{K��ҏ`�M^?�h�a�V�H�ɫ��L�B���L��n�f43���e��W��j$(x�ϪKt��jY[[_��g���?㭷���^d0[��Ї1�mz9�|M��o��6$�	�j5	*�yA�IAK j��VMKzYBBM�����{M���h�x<��"��)%���o��L��	�����Ŷ��Q�:j�b(������ҖI����>��3�dhS�w�'Nhz��"3*��*���
�_}�w�{���?���H�<9;"����$�hԱ85�j��䬬�W��!��S;��!N�<'IH�i;���j;)"��F�,b�X]"Ԏ�p���e��c4s��u�@ӵ�4��Ӷ��rfR{ �,�X_��/��������ˬ�.3�kO��M�����)K�HI/�hK6IN�(/x7����E#4J������t�Ę�m�8}�SZM���������j��V�9���ͽ{w���g�uzo�La���L��˄��4����G��nj�+�w&����y������e~���y�ݷY\]��5���OVSj�.A�fږ��vI��$��t�RSt6�ۉ ��ti)Y��>Z:F�.�(!���4�9G-)"ܻ{���vv�Կ��KJ$BA����+z�(�5���Z�]�9����~�2���/�t�++�t�#��D�Lr�4�8JDZ4`0f|�$���(�W��p�3�P)��f))��4`�rIqG#�q���Jۮ�|93XXbiy���U�77���f4�u�Kj����-Zr� ?��{�q���*��ږ6j��c*�,%��2U(R_O��2�3+>���}�{\��1��z1d���AK*ɻ�f�bz�b���*.���?�9o��:ϟ9Ml�" ��JPsK�� Y#��zA�$|P�eP/2���U5���ʬ���Vh�T'	A�/^�r6�C0�����I+~
�x���iY>��\׬�l*����sX�1I���^}�~��_�޻�q�� j�lp'~J�!�y0*�JRU,T�E�y�XU]WJ(]��d���n%>#�[��
���*���
$ZD!����h4b{{����k�wh�F����g~0Eq�`�g���I�������@fiq��.��{��;o����	�J`EOU�Q�7�.'$F����S��*�sT����0dXY�5�Z�w8�}0�P�ҹ��6��k*`�e	��-��� @�O�������;�j��&��S�:�܏7���� �,��V��y���y��wx��WYZZ"T��$�RK����">i埔�.��Y,������2�����T�Gj|�.�����!�R�6Y��4I5cͥ-uj.�|����+���>��}���[b�Bp�|{>��V/Kz�л��' Yc%VWW�K�q��>�Tj�o�JE��]t����>�-�����P��53�@&��b1�i�|��)�V|������%�VV�RҴ�l�V�#e���2�p��
T�pUE]�T����O�.�@!0��t��1G� Q�Gf\*�I�i�Kjep.�	8�i�{�4����aK2B�?� ����j1��<w����:?���8��q�ὕ%�Jtɥ�C\BL��.P�@U9�P�+=6�?�L�^�%��ԗl��!X�^�`��]�R��9�i*NX[Yf2�0i&ܾ{��x�h��s��b�u�Q�e����fم�۔i&Ts�����A��0����w��ͷ�䕗_�5�!��X4��0o%�$�)�G�*��� UE�UU�&��O��p-�w����j)I"��i���
j_i�apԡfgw�ݝ�ww՚ ����9�<��b�"�����3���;���[�9�<�j�m�bc�_j�9X!suJE��"��*�:�^*r�����y'�.�w*z�����ě���f�Լ��f�/����d2aoo�k׮i%���jjb/T\�A�h2�Q�T!�ɀET��sj�5"�_�<'��x��KA%�G'�?�!���������2Ο���~�7�x�Sg�cXy���DGLB����,�3�
���i��*�8�,V��e"�G��8����,(3�	ńDHA�%kc�iu�]α0X ���m�^��M�-�?�&r�wY>�y(�X��w0\X���K���������༣K��(s��'�9�Z�!)��
!x*c�!T��,��n;%������|�u��yV�@@M�UmDM�C�j�sܸ~���v�v���0�DZ�0���?on���vj�y��@XY]���s��_��+/����Ժ$�jS)3�Y��"��Ԧ�ׄJ��8o��e�����D���OT���L�)��I����	"�%�@��������;w��N� a��Oo�U�7<�LXZZ��W^���������Eg-����ϠՕ �\E%�|�z��o�͚$I���O��="2��:��{gfgA�$��b� �|�'�P�
^�_��� �%(�����L_U�]}םUyq�����S������:z����ڻ*##<���TMU?�����$�����?d�X��pvv� xs&�x�)�z�Pa�3<�j��~H	���>Ĩc�4�kE�j��-�}�s�����ދ����,���P�~�D�ڰ�*sm9ceyW�^�O�lmm�׫182bF3�:@Q**�\�|��=��~4��d1��uJ �d*�'�W�C�N�nT�W�6#G>|'���e�;�N����2n޼�7n���k���� ��?�F��D�a(C��޺��߸���Mx�ؿB�񞞴�C۶Ш�v�ē��
ۇI@�<�s�9+���e�N ���L�j*�l
��@������~oݸ�nA�������M�ͫ­�rB�6�/-��[7��6�n]C�[CE��`�InK����T��*�ޡ�֨\ž��Y�!G�/bF��u
�����Py�Z �*T�"jyr�r0GV��t:ذ�{+�+p�#6����"���X�/akk��6��n���"�����B�@�z=��u�� `��A��!t�.5?��&�V0�$�I@�j'��*nd$$x�I8���= դ��p8@����������%67��r�������(&�ֺ{�,���]�O)*}F���&�!��@UU�reׯ_ō�QU5����@R����1��Ҍ��B�� ��Ϝ��3��xD9O�x�9����9xWù�&g��2�'B&��e)9	�������*n\��w�~�^�)^˗�h���(heL\p�v�X[_��޺�n��V2`,HSƚ�[��H�-2��|dP�Cac�`<'�ۑ�f%�(*�{	��1`Ϩ�ȑ�� 2�״�����❷�fiEݥ���pVV:�$���U\�~W�����`�Dh�l��d�ɚ�[��ɂ�{��� ��R�:b��D���x�3�eQB�mE$�@��<*$�f��٘4f�4�E�c�&8�����������Rw�S�[殗�}lnn�'?�)6�\��)�k�mVDM@��D�T+���^� )�����ٱc�afˁl�GP�<��Ъ�K���:sNШhS�p<F5�76��O������.#�,��}��E�>�B�����?$��ܕ���D�&x_��_7p��Mlmm"��h��6�	Pe�d6E�;�P	j�0'$H��y$���2�rΠ]mWn�m�o
>��=j�A��d0p����#DH���ST���������N�Fߙs�[��)�kW���ͷqu�*wԚ��Yh�$�;��Ρ��
���b������4�l�x.X
Vc�6_yv��v�D����rK%���UEPK?���굫�v;�y�܄XN�YRE�]������ʕ�|�&�����ap|��r�-	7jh���z��j_yh��"���
V��-!`U���]T! t��h���^�+�Uؽ&1�[��֭����obyyy�[��W�_ZµkW����670��Q!B��i��=m���k�ePe[@��~�w�X���<�JRB�᥶�4F\�s�@h�#ʤ�P��~�:�\����2\pF�h��e�XD�+�	Vg6E��0�l���Z����;80������o��k׮��Yb��1��Ms�N�=CT�\_��S'�Ɍ�φқ^	�$��L4n��v
����BźF��R[cM(NP���>�67�����β)�i̗U "	b;���2�]����5TU���ڿ[h�HN�4CC@�T�F�+n�<��Oż`f���8�P�
Uͼ���ez��JY�"�Ή���⭷����U�m���@@�pi��з�G�;�oݸ����X[[ ��Bk�N=} PxH&�\����	�\�Ɂ]BF)dEm��U�����Ԩ|q���~y�"���P�F#Խ.6��p��5��,�S����-� ��*��}����5H��M�v�ӥ�`���XY[����3�c�SCI��(AC�/!xtji��<�.0t�bZ��e�U]c}c�k��//s52�Q.���>W����G-.؁I0�BO�����+W�����=�{�L�'ÅD\:Sj w��{W��/'��ؕ8^Ȝ��<�B[�˪g�B	H��|��Α$�Wb眔��rX�����J��Y����w� ��r�k+x��[XYYAU2�̼���rރ��ڣ����<���D)�9kT/gc#�z���C�QU,9Ј�� ������t�����:��o���S6g��`H��F���u]c��U\�vW�Ȍ��z;
���t�<$AQU�� ��Dѿ�u.2��A�
Ups�P���H�e�s�������W�3�4�oZ�Jgi���677���Q;�@�p����̆ �v�ޑ�)T�g=����Pl�qqO_�,Q� �:��s&�L���S@����s�����
66V�+4�5�`[�e��k��<)svVL��!���aum��+�<@�h�!�EP{��T.p�ڳ��%&
��s�̊��N���Z��9�`N=��lы�����;5�������n��l��7*��P�a�P����w����
A"Ÿ��%�L �P�3P�sF�7;��!�OR\V��� U�N��
.;$�ȉ�� mvL�,]Z������*��TV�ɵs�)�_H嫪���&�^��kW��)��������99k �B���!Y`s�5�N�ö ��F�ׅX�X�0=�w��pdpX�/ciy	KKK,�y��;W��ۺ�����k[װ���P���5Â��~�ZR�&^=7I�fv{o�BՌ�MPw*86�%J4�foz�y�8Gz�����:�a�A���b�&?�%����@U��P���*���h[��mV��en3�^�+.Ɏ�' c{qL��XfA@�cH0���>����0�� -��Kސ�I�������o�c��'���	卉��'��
�B�����*�N���� '��'&\���4B�����E`,���|�Q�
)!��'D"�3�Ȭ	�J+�$������p��ut{V��l����I�(�4!�|F�~���误���aژDUĜi����Mr�r�y@��ܻ̟2�Q���Iv���d9�l&�$t��7RB%B�$�re+++��z����r�u:XZ���!猦!ZYr�Q�UJ��mAe�T� ��s�so~��~�se�$�$�L��Y[��49Y=�:�l�_���˽*���\JΝv�������W?�{.�7��2//�,9q�QU��.�u_��|��9zv�ܜ�9x����AF���=��\��;'��f��ُ'�� 	�E����z�"��'p�/��}�˫�-��2��!��sF^4�t��*\`��R��~��*x�0�>�<Nr����t�V{y�tgF������b�$���"�a��G�!�t� 7+$�r�%n:5���"����2�8җ�)yۄtЭkt�

��Z.�:5g:C���޻c��|���"`�M�8-,e����xe�:���s�²)�e,�zXZZbs��/~m)�0��:5VVV���J�3e���ɠxȞ�*��]e�4��=�2�_i.��y압\���� �^��t�Cݭ������̐���e^�u���C����s��[��THS]�8�dT�N�_ʝ-�ボg�s6��`�J!sh3Z������n��)���-�rW6	�3�:yOɽn��/}�]��R�b�i汪B������J�]�_���d��(-��Щ;��GΊ��
��E�I��_��E����.:���@��s�ȬYsΑ�G�;�E���db�����|v�U�H�+D	)g@�*�h��ZC�v񵔾�v�7|@�a�d�<b$�+y�Ä"G� � �Cs��lN�e�Ϳ���e>"�3眐T�Y�
��
�Zfqz�(�qh�gU�F��Lxlϟ����sH ��$"��.�K}�����"xG${�}����;����RH%�~��{.�E�>���^�Pi�5|$���Bٷ�{�QI��K��u�zP_�A�-���٣��r�p
 U�)�*!匇8R����'"B`C<1j�.�>7�Ϡg��≭�vu�3��L!�5�^�M�2i�7i�]
*�L�`_�p/s9�}s�uz#�k@3D<�d�.���rb=�#�yyj��A�Pt�O;!}�X�x�!Ig|�32{J};e�I��5g�9���bm�JSj��t��1g����<b%F*�� ^^�a$��Ia���Y�<[�1�-H�١C32<\`��Bm�0�e���t�^v<�6;f
�.+[�	�{WD���\C9<��9�r56���]����/�<�n�J`�&��9�^U7�K��Ō(�˅�^fr��uq�c/�=/�!-�{N潋D�5�1�^$�jt����Ρr�x�s��?��#����BM�؉ɑ��
�3���Su�����W�bksK�.���Ba�]���3;�r���)�7!�;�dk)�爖�ZJ�ą"
��#�E�P.��ˈ �DR6�v���Y	"C,�Lc��d6��@�7��x^��;O}�����%6;�����)L��g���iX�y9�����#��SGL��N�:�0����=Ng%�1}!}	qENE��/�~$�U����"�+��y\7HS>W�&D�۵�{n0](�}$��#��m�G�t��C]��d
��k/!�!Ҹ[uP��Y��mD�;r͒9�քL�0]'(�P�3��"��<�~�����,`b�P�K�e�1����Y�����,G/c	����,\�����8Al�;���q�w�ӟ����O����nw	�W�N��(/�G� #V���:�d&)�	P�BcDBDL�|���}������KY���:V��5��&'dIH��ڶ�L�5Q�á�׋vҋ��U�����Jƕl�0)�8c��*�LP҆%^L�;Bcz~,^g<�r����Y�"爜[��P1!�mL���~�΁�_T�q����9l�S���4)r[�`|�<f�=�:D����>_�+i�ONC�)ٳ�5�ɰ5=8Қ�����z|sBCL��4�Ft�a �F��<���LD�q��s��� ��g�W����q�=9Cs"(M ��KM�M V���@L	)��֐�w+���7ϏǏ�H��D��2ڶ���*���#���?�������+�������?�s�O��?�ͷ�B�ӵN�7���2W�4ve�M%;��Ӥ�.d؇-����8+�?���;�<�\�J��H�Ч*i����sc�����2�P�#
��I�?�=�p�[�ǰ�LK &�C���_ ��n�Ӕk�������˥� �i�T�mT3����|�3�E��*��Xa2�����y�V�˼au
u� ��@��/�3�����(��V�s���$
�[" Ɉ���x��z����I=�őJ��e��4y�u�#g�!�� p0��B�nc��J�9Hd.��8e�K���H�/����c}}?�����_��'�?������~��g�?���!�}�],�{�|�#ѹ�����0���Z�v��{H�Jn��Bw�b��70�4^�FE2�rcO����*hLs6�S.CJ�vơ~×(�I6��<;#����p�Q�=�ox	��3�(�N Y�����������,��ј���&JT'f�U�T�g7[ك�"�e�^nv�����}��qiQ�����"H�Q���s��EG1�`�«׬H)B-o�j=�){�xkG_���̈\x��(���c��ǋ��}��c(Z�"�
���Zf��b�Y�q�p 2�.{/X__�;ﾃ���C����ظ���J�G��?���ϰ�[:���}��I�u~g8���l�A!��U�$��)�L0Y�b�M�S	�#��$h�gϨSIb��qٵ����g�m���xL��SO�j��t�{�������rb?g*�ג�Ϭcݙ�`�x���"tἢqrzb
��3Chs�ޜ��X�5�Q�u�Y��z1
z*T��@��r�8�\�������?�I���֙���U*�K��iD����y���\���`x�*���U����\��6A�[,�AT��	�\��Zm�S����/b%Rbuƥ���3�l� 8I��}l�fk���y��嬜��ZT����B�Bo'D��#Aж-b�h�!x��ˬu�;��C8J SD�DG#�UoQ�z%KՃ�p�7@�!�$Ψ���!�W��"�9L9��ccF��4�A�5���P�h[��M�0�Z�c�	qȀ��A�f���CB��L>[c��tD�c���m��Q�ų/r��\�i�hitn=�x
`��R%���Mra xR ����ϖ��$[��X�_{�c��s�|��	�������Ź��v���e�Y,�!6�Rb�N�����'� ��8W2h`0�m�ϥF^Of֝ ���3NNN�����v�b�P��d����%<G?w~���e��I�͊ b�/�Z��g(�{����D����f ���3B��r��,�a������y8�h<���	NO���);xqh������ m۾)���H��s���p0ĸm��1Ө%S4O.Y�!�4�)8��P@pX�2GV49�M-ڦEj�S r��D�MsF+
��b8�m�899�h<�����oJaM�Kj,B�	�m����-ZDh�� G KB���آ�	���鉖����ˎg6�o	 '��-���Ƅ�d�����Q9bl� �h���bJ�B��d��H��H���PI:k��R�x<Ƹ�M-�8���$�Hf'��*�$�u��1221��s�����8rJ�P�ܜ�1[�7( X*���K	P�#588:���)�����ߌ�� �1F�cg�i*�t�졚�Ѥ���8���)@�D����RF!���Qm~�猪R�"�	ml!�>���+�Xr�X�2S�b0`4<E	$bMЙ�Q�y�{�:Q1�j�)���;�����c�F�� Z�pp���m|�ŗ@��MT�<2�ض89=E31�#bA5�)I�dֻB���hsF�K,!��x-z��"N�SF�	16HP��쐁 �+����S[��J������$��J��NR��-FcS8�l���ȄU����&D����)c��w*�8�b�Hm��&�<T��+�i�0�p|r�6FhR֟:2�Lc��ฬp�xG����ǈ��npN9�d���Sh�hr��xqI��\ ��Q���;"Rl1�p	p�QU����FP��8<<���	F�t�~�"*�1����{hr4:�)hNDH�X����S"g�ِ�cw�/��>D!�e�Uf �&$>��1מ\��9TRa4���'��M��Ҥ�܏�bYl8gD��9)6��JG��������_�����������?�;�������������p:̴��~���p�9^��iqr|�gϞ���rnB�:M-bn� ��@����H�����vNӭ�9'��2bvsf}&4Qѫ��zXx>!;%Y�:�!�����w��c3����ʙjG����O?���!Ʊe�vP*O L%x�1s$��EkxRZ�M'�{-�*R�&bԶȩAv
W�z�<;5�S�V�x������b< d������)�6u*�m���<{���{L;�LE������|��������~=c"߰�5Rf'�6N�O>��R
�@[u�����N��0��إ^S|vM�����̳��ȇ�]p
�!�Q�x�Edc�<eQ�ȅ�}�Ae�NBBJ-�B��W���I�;���6�8>�����5��������$H�+�0�d�)>��C��W��_��_�?��	���=|���8:8D۴�������<�X�Gezz�gϞaw1):����,\�N�
릑�c � ���R���Z���k3�NQF�C�gl�
��*2Rj�X)L���`
�&58q����CN��?eXyC2	}hc���!?z��� )�	ǦZ�mIɪ��'k�Zݷ���̶N���{�ۜ�1�HwB�2r�"��4&��|�:���U�U1�899����f<Y�lyj����hb���]���a�N���nZ�č0���r>z1
�2����\�;&v�Ρ`�	'�&e�PWLQ���c�t^)r�C��cF\�s�2j驜Y~w:��t�h�y�dv�9k!��L��Mf!T�)����5�(Լ|���� V��[@h����� �����{8<8Df�՗��Lo��4����L��)E����7��~�˿�_��_��o�Ⴧ��g�鉞��[�\�/��U��Z��B�-�!���h��Ϟaog����K]6���yԵ���jB+-b.�cC4�	�x�8n[�J�n�`ںl��CĚU����DT2��B��뼑�����!��qtr��x��pT��U�#� ;���1���#���P�k��1D ��i��-Y���dc�a�y�n�\����䭡'�^X�}@v�#���F�$(�g�Pf�A�dAeqh�Ŏ��&%��P�.q���e&)������F��cww��ħlC�0��r�� ��a��~�!r�J~n�M7ksG��H��FG@��K4��v3٘��N ���
��+X�?1�1���9��:k��>29��C��4��!NOO��<�7�8�
d'�@�B�Ɉ�yP2Ky�^��d�q�g:3v�gEx�b���ץ��L�Fnm�ǽ�섢��h���cq�z��G�+��'��[�712�ГR�!�ـ(�e�Xs�Y�	m�hڈ�#�8��	Μ�;$Zvb�a�Ҥ�� ��?K�677���!<4&�6"Ó)j�	9;��́%������������B��eP٢,a��(/�#�ۈԴL���2��&"���{�qtr���|��>��o�����P��F�k��������BV0U��.67ֱ��I���H�wAO	h��*�B��ROΔwQZ�Ɖ$�_����ZZ��$2֞�b8"�Gllf��޳u���p�h��p�/������ܻ�����FE���Ǚ�r
I����YN�l����L��ﾃ*�Hm���Ы8��EA�
r�U85��T�g��y)�iqלkÆH��m"2��;E�pgAqЩ{�����}�?�>���	�0$�{м��׭���!'��F*��
�N�+��v�����4!���  fЫVE2�cQ �昔�F���e�����/�ɠ�\U��q۶�[h�D�B�s���8F����Ɲ;wp���O�� �FfF_(F�0���Ẉ_]Y�&)�E�[_8�g&�+Ph�T�m�"�C���Ǣ��Mw�"�RJhF#��aow��{��1��U@�
����gdo]VrD��� �hb�.QS�syE?�M���Ϭ�R�kۢm#bc�H��D8�+
�E�N
@Dʊ��	��������y�	���|yU?%��2��*��������O����&5H9�OP����^'�O�A�cօF@�)�� �q2��*�*w5���q��f�y�N���X
#@��bPQ���<���Fá�F��%i���Ή�\ �(��Ay
���88<����wѶc�NՄ�]�g��9cİm�6��]�u�
��ف�s��(��n�q�)���� F
���M����)�����c<����`@D2dƥ$��#37:/:ʨ��Z��vvvp��}���Ac�)�H@.�����MMN��"�mn�Sd.188�����R���l�UA����Pw���|(o�I�"p�H.�mZ����ރ�����`0�3�����sR��e����]��IE�Iz0�LȳLȭ�;�"ԑ�)h�k	!����!������m��#$ ��F�d@�>3�瑓C��c�
�������-4�%9��^��X�\|���4�E;c�4h��Ɇ��)/��ܖ*�z�pzz���]loo�y��t�R�DA�U���.�iZ���x����p��d4J/�̽Yq����	�آGhˍB��:��1�{�6�.��"
EL-FM�4O)#�F�k`�S5��&��� ��������p8�.*db`��0���uic���v�=���.ƣ�{=TU��R�!��0�D��(�<n0J	)6h����f�=�3����p�(�H�96�ű�'n�ٓx�	��ۀ`�&��p�O�`g�f��g�q�&�/w(�-;uDD���G���èiX���&�F��n=�M;�x� �ّD#�آ�l�1f�z���ֶ
�VO����Mc4�͸e�Jt���mF3�K���k��/������`%�����Q�����Mk������Kџ_��7����q�����e��AТ��a� e.�N��R��Ս�,-!tk gd'��"��8`XVQk$�`��(n���P8/mC���B����eĶE3�'4hx����@	��\t{KHM���]|�����Oq��7 Á�%9�sM�J�r#�М++��C���u�յ\�~�WV��t0َS�ͱ�� )�,t�)f;/Dz��4V.�PY��K$�匤�R�QB��HF!ʒ��+ᦢ�������c|��g��Ï��������V� ΣE�j��������f�c�*�'���VWV����Ԍ�T�UC��V:�6�R$y��88)]}��OtƢ��I3T�!�6B���FV�$�s���^<:��z<�y�O���ݻ�����P5��83�&���ߙ����2���5�F�5@Ț�ue��[���&h�Y����#H�H�j0�n��MD��-�)f0�d%�V��`�/6c4�E�-	41nQ»���q�l`j��?x�O��ů�{�{{�F,�̕2Z��9_fG� 3��sgKm�s���R��]��ՋA靐qS��D��"T|Ua}}K�KXYZE����*��3h�̃�"� d�DT$e�6T�Κ�
��43�̛*����h�zH��>�P8�&�"�B��Gfn3T8��Ⴧ��o����
����m����& ���e'C��	�R PF�@SFTv���z��������fo������A�)�����i�S�R
�K�bNZ� )�z�����ض-�� G�8�7�`#���T��)!�����ŭ[���g�����MV�Yқ7�b
P 8��C��^����VWWQw{�bݫ��:nE�iE�rt@h���H�Zn��H
�\��ș �&F�qBV�hE@��p#����:�{��Α��S|����s�|��8��g��B��������A��T�oq~zFۈ地�����e\�r�3�NXX��ܠ��K#T�
1�jND�j����85/��,D⃜3rj�c�8F�'��86��р@�-N�TP� k�x��ӻ���ݻ�{�.F�Ѥ�������E�x�~o岆S����d���z4�~ȋ��,8�F�c����FQ�읠�~�����6��5"fE%@�Ye�p/tb��3�6#�EL
�ڜ��1%�ȼjT��1&�Ѧ�mj�ÄQnP�#E���.C#w� ='O�>�_~����=<z�ǧ���Z1/7�������u�0T��C6��IM�&l^����
��]�mC��0���ن,)�DQ���mJl��"bJ,i[��h3�)m��6�"��q;�p\����:1��`ra#2����m����}�1��<z��`��
�F�����'������ו-��n���\�~
�h�n1C��X9���Mf�G{nY3rL����m��;2�cLh���9���6(J/'�)ݺN��0���Sܺu�|�	�߿�62�0��Ύ��5|�猦��	n~�$.�Z8Z h�1:UU������u�
�m���2A�d�ҼŖi���-�w�@Nh��Z��#��9"5djR���Im��Z�9�e�cJ��Z�9 M����x���|��G���]<y�*� �5!���l^�7��������1����p�236���ˈ�8�Hm��`��m�7o��N��^��  �w�"����"/�FYk��d
JیF�imי2��cn�(r1ID�%@�G%֭��$�"�G''��O��߼�/����GpBf[6[�`"L�r� ��Y~�x�`���m1qec�+�غ�i���qۢv�P�^��i2\��K�%��EE2J��
$�~���3KB;�m2��W�Ly��V��̏�WC$c4��۷q��m|����Hz0����E�iÉ3!}�=�1c88��u]a����>zK5󵎆3[��0��T�YA<�@�H1"�d���#�I[4-�d/�!R�{�9 `�fj�T\@��������+����߻���#n2�\�y�Y�f�E1d��u�ED~���`�e��<x��`}m���V7 ��<�0�"���"�$'8/@�P��K����uc<�h5��Ao��A� ���՚l�C�W{��V���2�s���Ç~�;�o������H� ��ԅ3�,���[��p��B/>�;,��! pܵ�q�4�U�����R��E�S�OU!j��u� Rf����9���#2���";�Ė���"	A�Z?�LĞ�ܙ�J�"p:��/?ǭ;���'�����a3F����~�D�����߫'�`�+  *�|�HJ���>z��VVQ�k���j�r�k+3�: +��@�u����OK̄�m!9��	����ba�S hsD�+dI8<:����G�/����'��d��6I�Y��g14x�7fX{4n<k)��˨�=�./s����h9ayP�g���-b2�5�����m	oVd������乆 >�6� ��`0�_~�;�?��;�����ј��B�G`�s����1����2��Ԉy���5j��q0i1��KTz��^>p�$�P����wǁ$:�!���<QkJFx�\jJ
$��C��h:����i
a)Z���IMk�b�����l�}�9~������_aww�!`e�`�T�в$�ϸ�R��D~4�S��^tP=O�\��PLM �laU��+�//ceu��ќ��q136=�'̧��1��2!2���t�F��-��=w��WP鷒t����@�&����x8³������O>�W_}��6�6�ɗ��/��N��ɒ�A��P�%�p����1����
VWW����E�֏
(��C%B3�t)E 3̭ �e���z�jBۖ�"c4�苂��j@ �LP�	���N@��C3����������[x��1N��3����jyNE0��k�On����n��K���D�� �A�)"'ˡ;7Ť�XGK�jBL,��9�c��#��A�㉃� '�IeF�9Y���y��a������x���������'�Xzn UJ9ʋ'׫���un���YA�	��o�qCb�d4���`ei׮\E3��wI�'� �xT��{G(7�� �� ȱA�	���9$��p���I�!�p��s��p�������1~��{�� �0[[F�wV�(�@�G�yV����@{(Vi�H�:thc˲�ѐ�Q��S��uѩk8���� ��`r�	��Z��	E"��^��f"K5��#��2h8Cpp���t�/����~���x����!=\�F�T�e^$�7�(�f��8�0�� P����4�S�ѭ��6��%][�]]J�EB:��EX`���Ώ���F�F@:����k�n��oy�����̝s�y.F�	N�lp]�|Q����@r!��Ut5{���3q�<	��:����gNgx��y��!��V����Y�5�������9��_p�V��?{rU�)�W�!s���U�&��,"d^���+xB+���ڦ�VV�\�l��r�;��.�WYu@';m��Ap}��V��+F�g�M�
t�Vĉ�����jf��7�	s�
�Φʻ��*6GM�o�Yv�1����&�K����d3|�4/�D�t����m�囑p>P�k/���GF^���8P�I�#��sO �*]�B��ﭿ���/m���L�G������I>�T�Њ�\P��+�eF� B��	Yc�W��Sgp#�k�NT^ô������//9^�g%9�CWֈ��
u�v̖�c!m�ϛ����;�}���g����~H��S������x���a��(� T�p�x�^�����8���8���kg������6��$�VuC�S�;����p�֟e+t��F8����b�ؔW\M_����1��fqm��EF��@�f�A��B+c������ʾ ���~�_>�C]
ƴ�9ګD��!���a�z_~��S������D&��	�-��؇���gf	V6�������P��=��C*�\��F��A��<C9��(�J!2�A�I��=�ؓ�jb��L%�o�4�	lr���e�/-�	�$�_���8��m���x�Y�:�{ݷr@6(��u6��b��wԙ:r�-�]���W�L5t�N(��vR�V������Y�����<{`bs��\r�@Q�	n���4��VT͋�]� l�k�VQv
p�#F���={t<�D�ٸb�Y{zD	��*�NZ�(�6�M	&���Ft�\��O�}F����I+�t�������t�p�B��Ĭ ��ܽ.PZ!~�z7E�ͯ�{�A�S� m?,8���I{>�+�|�?n��Ev��F���q�-��t~]x��'����W��.�d�[�P�O3e��3���h��M��f���F��;M�S/z��A����~å��~۳�"���2�|#���B�wFr�W�@���g��4������\����D8z�P�����A��L}���z�ޠ0���✍��'�W|a/��=*6�:w�4�R�o�7?*S�����Bo�!��'Lr:�=mlciY��L
�Ñ]�����BY\��ּ���4V������!O�b'�08�<B�jͷ�7���괐q�%D6[w�u�#oXG,-5���ݘ-�{{��.�$S<Z������Hi��=s��5}�	X������
�p���OZ��7��i�2�膓�9iu��U�(��Mlp�ax�.h2�}������t��c�Ryߒ���>m�~���G�2�M%e��W�C]�i�:c�5u��	�4�D��a���7UI��R�"���9�MtR�e#��>���j�s�yT��\)4ǅ��	��ێ�4�X���ہ䔇g����b^�ņ}�
<�_���.({W���8����fCITh�'
��懡H {kwEIO�j�yd�s�*��]}���B�ف�P��J��)T�R�͐���[����F�b8�PLQ����'TU�q�'������w��1c :�6������E��F��,�ߏf��0 x�z	�C�E�@�J�(�@ܺ��f��G'GI��g��4k=�����8��dr�:��.ޱ���z6�$�z�$�/,H2�g��ǘ �(ÉeW3�pz�Q����`�������m��(�}k.aC�A�E�7-����o�����S�Q�I���`�v����A������S��rr��Z�@����&CKE���c)$$9�sʦ$�ܔ�נ�h'QK�/�ĸN4�&"r��i��
����`j���Σ���⯎��YaX����=V��VWW�%>ڄq�>�3����\�sfC�����'��v�=E���:���?��T�f� �����G*��^u����;y��{R���U�P���r�I���Ξ(�\�w�]��8��9�f��Q����&B9��)�)O��l�֎���aw��,,"�󙀩k�z�*S��|��۸�����tѭne ��ǿ �ճa/�TL��1��1�~_c��΄'Mi�W|C��E��������7�a��f���0�b�܄I�_������`���|I'��G*���	�GZ./G;�{��k� )?���VJP}swvX�x�)�i���1Z�dB��՘�>��X����v>�����7X�r���>Ùs�7�������m�Ϙ_��bx��м����ВN m�wR����^�,:%��⼸k�����;3"�|��ϼS��a{:�(��G!�xH0m�!����� ��w|w�{���,D��K�P�Lee��x���G��i��O��-��+����m�M҈ˬ���ed�~��~���(�I�9L#K� ͣC�>CuEG��fgZz2&H�P�.L'�����j�ҿg(Yb���U*�I|��v�=g�Yג�1{,�rWF-�]І��bO]z&H���i[[?2�&�U@�.W;��!��N% l��i���c�w�jvv����;΂�)�'��qN��&oKǪX�A�7���6i���j����zm��~J\{��+�龛���f>��lJ2��9K*���+����:���)��7&�WT�_�|=%|�H}�{؋�_�X0�o%z���Yp�L�,:����88��/����J�~^�E020���6���XȢC�Ͱ�;uHδC�멁�J��!��A���(נ0�U�����@���� ���q��,5�sܼ�Zz��n����n8^<,��/%����E�E&���.,d}>��}\l��#$���9I�.��F�X6棠��\��C����z��H�m�IV�~$�`?�q�x�
G ��	i�BŁ`)�Y��z��8&ps�H��$���G03���'�x\�KJ#'���;��߀�2�]�Ͼ�y�$t�u�ݝ��>��R�Pļ��
z(����~I��hbA��A	�x���*D�1(��v��-0Z/I������R})!`�7Ҷ^z#,|�x�o��z�/��s�~|\�(aS�p�uƦ;�r�E�Iݠ�������f��"�{OW��e���8E���@�a�E�K�������_�_�^���>Y�h�v��à�^j�J��ݷR��3��:Q�XM߮��=��4�}+ �kp��ן;�s??iq4�9T���`�$�b> k�Xm���0�`�<��D���k�ꢊ����֥^�c�E���Ɲ\<^)�B�]=a֤�ק�c�D�-3F��cLq��=���%Cd��+2n�JKk�O_�㧭xpȮ}��	�Z�[����Ň�m��B� X�4�S�
�B'y��!��Ɗ/ꡤb�ꋯ�j�4�#�ݛq�G@�&���!�x���?���������)�����3`=Q�:�}��Uȟ���uǼ�;��y�q\�ƞ�2�<��<L��o����f��K�"U2��H"�wޣ�xD��P�P�����Q�u_]i���~#���G(Z�&�gN�vg��_�N�.�f��i<9���p)6u�Cu���R�S�)c�7j~��Rǎ{~��oĶe��������=Nc�sv��x�]h��Yu�Z���Q�=f�E��c�%��=��?�b�++tz�qᕲ���W������<���h���R+��k
���6�A��B�pN�s�)�d��1�D8;W���+Xu�����ѹ�ٌ;1z"§���8�;t��t�m]�F�32Z����:b�����̔�8?�}[n=�:7W�|Z�1�3<,$�B�A٬RZ����{-|{Ǐ��4�D2n���$�s��p���x���@�N�������p�Ԅ�B�L����[S���㓌*WX^%[yy���0ɗ67��J��ׄ*�,H�5�mo(�����'v��-&^�b|lLA���Ug��W�w2gO���M�#���$���՞�.�lў�I$�8�<���j=��P�txH7A��E 
�Y���|՚;wl��T���U7A�23ujΛ��ퟗ��gޜ�dq�FH���9 =��C��?|�	�0^M��P���ɉ�������w�8Y��t��`��J>2�d"��_�2C�Zo1o	��CY�R�B"�#����͵!e����l�s�5�K��ǒC��T��Y�Hw���6L�������l��N����qg����r<+� �5}O�K.�D�d'Hj�'<���h��9�j���?}����"}� ���yh�C��f��蹺z��o�n��"��8�{G������>�l�m��
�1 m�<S_�vDyU���ZY�mc��r#�����(v���C{\��+Ua��98颎��s��gYZ���C�����b�𜾺"X&�ז�
K�pݧ7�|��'�p˽�i��������-� �_�5R��K�����Ĩ|�Eq�\Զ+w|q��Ȉ���G���~�қ��	~��{Kj9����c��Y������>i\�ӥt�̓���(T���K�Zh�9_�w��PS�w0c�蜕�X1�Y�X�u>GN\(�h�L�=��|l�
}vz��d�,�u!6�CK�I8�e������u�J�u��ۆ�y3����z �_�
Hz��`���t�p��X���J�iw��F=)*�����.�X��������ܧ���<��4��I����R��&��5��G�Sj��!�'�nD-��^=�h�^�� n�4wߪ�f�|m�"i��"2pcqV�!���l�y�t~qQy-�nY����N��0��{���ʠ��m��d�@�����[	��d���4݋#���^,F�[K�!������X亱����Tre��E�$�i�]��=����SaN0nzk��t�����`8��\ϧW��/<�*�w婫wb�X�qh���t��0��i�Qނ޿x�����wI�/4x(�~�X6��T&Q�ʩ98����/��A�х���^�wBb-0���Dw�L�U�&�H��}�����@����i�T����0�Ef�~������.Ị9��Eʑ�!̀*�}"��O\�,��E�{l(�vG:l���u�͈�#�K�jq+*�}�Qlm���0*���`�te����<�P�PTc�j��+���7��8��^���8�Ivw� a|�d�!l�݇������؆�戎� ?�k�̈�i�h��DC���ix���{��݂���|Zg�E"W��H5�X�cK�U��a�J�e�d�OrO�K��~O;� �O�<��C`I�
�H:W�:�99ʜ�ϰ�1�����V �C,���S��zH�cg\��qͥ�3l�N9���j����*����������X��},�(s0���U���G�T>a�V�!�o�Q�8�ɇ��T���s��=>i�9F�&*��� �[��=���eZ����{ף7��j�D�������7��c?N���͈��46�l.R]��x
|-���;[����*��G%�`�?d������*����j�>K$Y��!(4+Ll8j�7ή����c_G���3*��A����	L�o$/5���I����/�Z�Ɵ	��ǃ(�
TC��
t����C�I+%'�\��e��B�ۢ�Җ~d8��6r|g{�?�S�OJ��G����v�����J�xB��n9r_!��#��Ъ��k�5満�$H-��*�*��� ˝��.�)�� ��y?�F��}�}M�k�;��O
GÀ�Y�@�"��<��5�p�G��7�DK��f�w{Ĝ� �}�����o�/݆;sb���jI�}�b�O�H]��.�k�G�������C��cʊը��2�yi��]�mט��MA��%��Fņ��z�X<D�w�=����$�����x����C���R�泗>
������^�=_�mNj��I�W�����lz��=�7MrP*�>����v��D�'Evϩܣ(�<��wpd팆��%���n3���Ti!k�a�>�����-��j����8������ٖ�AiO����.V�Y��Bo�:�-�!���'��+5*�M����vՏ4+�L�p:h�0aIo�C{�
M���R%!(�Y��6��X��ŘO��tL=V��6GMo����3�c����.��L��?�`C��%�M�fR�İ�y�Ѱa���#J�c�E�v����_>n��ⷕ�E>��H.�G�+0yH�:Rκt�|J�1�s���~Q��\���]�P�0^��!�lVut��j�&QLv�{-�c�}N�s�;�����d�?��w��EGnK$�[����A�JZ\�+�'!*����B����Iaɤ0���bHŻ-�Q�~ ���,��ݜ/�&uq̵=����)�aV�L������`3��~-�`��o��>���[�}KPu{KL�H�,^9��>��)�͸؊��{��<�A��V�����Q���j���}k����l,���� g�"=X�0�5�\��- �g%q8 �7XY#��fG��i�����0pi�}k�.����\i0�,gL�￈�5���$b��Y��j��Ӷ_��L���x��01d㽳��� +��2��bh�����:+����v�q�rw���A����ܓ��r�u⥠j��o�����(p����>=-ˏRIV���D�T��n_>w�t��r$����ײU~�D�Mv/����2�M�L�h��߽0�k�]␪`B�*�'���h�s���ͣ���\�Ꝝ������?��ZٙhE������2��-@"xʘq�˰a	2�?c��楩�BZ��ߣ��?�;)��.nE2����-�Ƥr��/I�8(:��b�<���\�d�l4��ie�m���,��+�S�[{�|����(����w_ fy�̀ԝ��TRh��pL0��7ĕ�W��v��Qp8W����h� �p���X_���)\�G��xXW�&��/����_v�mSq�C77r�9����o5�^*#�7����8=�M�(�W`��"�u�"�{��;q�
�����&��ˁ��h4־	۞�e���h/i�t�6R��Vn���daa�1ǽ}�3J7�����33�kd�<&uϿ�w��s����GDes�\�?�+XZ��jEXG3��0Y�t3.wp�0�#��8�'�$�����`��Jp���v�9�ǐ��)�%?V*�L����!4��Y�?4,e+��������������*�;;Ex�R����%�_ �	K8�T�Œ��a�4T���ƻ�G�O�:�ڢ����A����/Io�4�t��f���z�m��Z���3]O���C����x'����G\�i�Zz�7➐<���h��ڨ�����݅�ƭt�`�Dס �"3F�ʈv�xړtJ���BO�?]�]\�f�������H��J��_)����?gu�%�P�_�܍�>�����A�3��@T��e6MBAh�0i�Sr��~�T���WMz$�OS%�gIT�|%�o��Ti��Cp�w�I_	r7^ y��d��7�]���mw�Q���_�ƪ���V�DN�Z�Ý��~�s���m���e�����~�i�ۺ�����%����CT�qeGa�|Y����ͧ5�q��^f�D��W8�t*1��|V�L5�%���<m�a͠��Php�2�f/C[��Y�U��j>��k�c�SN��E�se�m:�ս�G����v����U�r������:J�������Y��~d��a�e�w�J��X��5��
7=��>���e	p�o�5<����<9�u�Lh���;f��H�������-!�Q�>��0��&�	�������p�������n�vh�,��r9�~�.�<���ɤvÖ	K#i���@]�:�o멝����Ju>���l>,�+c�.��V���B����H��Ί��|��"��F�3��&6�C�t��9ԕ��.v3��&�3;�K2�K�s������teZ�x\!"հ\,�N��ؕg�n/��&�m���c�F���Qx�*�|�I�÷A�,��/��{�{,�X�fM%皷v�k<s.����\�5�y�i��`e1���>�MNK('�4{���.��*;1�ا�k���5����3�С�VO8��V��9ea����oR%��n�q�����������7˶F�Ҵ��\O�ۈ�����G���[�~}���u�d�4�Y����ιd���^�v�\��Rj��2z>}�LE���Kc�;_9�u<�ѽ��_�̡s��d�N'H����: �ݐ����*�):t�K}��V�8����������+��Y�����[y�db��n��z-p�è���xWݪ(��ɋ)��,��*!�]��mM�O�ȹ�l�.��6�w@ �S�Q���4�PK   O��W��ܣ]a  �d  /   images/7cd0bce8-56da-40c7-a6ad-eff1f7eef46c.pngd�XS��7l�ҢAR��f�tw+�H0�V��!�2dt��t	�Ajtw�{�����^.v�p������Խs��U��q�p�ݻ�� /�y��}U�с��yɇ��}'M9�{��u`�JBE�޽��+SL`�Q^���=�����N�����(HKh�o�us7t�<��>�%{qޫ�G� ��AЕn�є�0��%�G�U�x��CZ�o�^�
+��o@G����@��'��
����ae=}������y�������+�M���uFɉ*<�,[�`d��͸���8��p���e({���;A&����p��"�i�L�@ �"�����c��E҉�3�3|���Cj,LG�R�T���Vk;�ETyb��S9*�*Z\��)Ŭ�Îg�<������u�uE�SE�G�ŚEa�
\�Ԣ:�����N}�s�K����_7.��Ԗ��7m{��=�Y�Uʛi�K��<�Lu,�q�x���f���~7o|O�3�]6��T�`i���x��
�8�+Q���k�r�f+��"�4�Dy3=L��J���Ϲ�]�^W�\v��\kR�k�i����,&Һ��M�f���:��ٷ�q|�}���~d}�bb
G �O7-�� h0���!��_��%&Z.�KuӴ_Gm���Y��t2F�a�5|��č�|?=�������U���S���~7m����0��m��tYBLTX�@��!�j�� �֏�n�l��0���Ꟍ+���t+���
���/����Mש N��⟠�oE��i`X���*��9sx�ӊ��{9�ob~����Q��V~'&����+mӽn�JS|C.�"_p���s0}_=r�@�	D��tF�������x������$��z��Sbܐ���2D����z�ݙs���}���\�Xd����f��ނ`���=$�����@�V��b�f>��u�D�����Ls�4t�,fo��]�࡙ӱ$F��
{R�(�H[�[��~�����o��*
y�Ϫ	��j�L�'�����2�A/
]V��OB2+mwdݧN���������x��p�5�D��tc�����:
9��u{�[�;k�*3r��}���ĺ{�k>�\{e�P7�)&�U�=��Tg%m2$�~scY�������ߧ��������x��_�d�ѡ�'Z���٧i��$��6�΁b!�5B9j���4�GJb��n��.��jv��D��1���9�[i8��B1y�}�|�-�����K�Q�N�(��C+�d �@�2��G�A5m��iX#����+�i���du�{T�v�iNg��eްǥ���c3�as 6Z�ƑjTG�L��L��!���gG�ġT(��n>�J��J��ߍЦ؜��ԫ{y�ӳ�-_�/Q?ޫ�ȆFoC�qr[��S�d�A�i׉�I�����P�✠�<X`�9E����f<������F���h�
�t�%��cTJ�)�{��3���3n��s�KB&I�D��X�<��ĘM�CSc��^�ק�N$�j}p��0$���nB��s/i��B�[(hX=�@�e�F/-�s�a���|�B���Ƃm��/��L��[.�����0��c����!t��O�ʗڬ3��C#lE-!T�c?'qq�s9+�
'e�{]��#.:~�x����f(�uAf;~�k5������Aq��n�:ڂ�@���и�ĺ��`q��s�YT_����HY� -q����/� iB^��3�V��.�v
x����`E=��@��Յ�ؖ��y����X����T�upE�6��_�9<�\"�,&��:&^p����,Z�d|�y�6h+��k�^R�%�d�|?ƯG���uk����i�Y
2��9������r�N�Y�k�_g��~�?.Ij�`�0�Q`{�_YurB��UV�م��6��Ԕ��c����1��waW#��ʡ�K���,*���u�Do���򩴻�M�ւ"�r5'���[�UUc�u��M���:��1|d���,Ƒ��~���"�����ǆ�{�(ry���\�/	_�p4u�ŹH�����A��,���x�l��oM"�9���f�Ё�k3��g�O��y�is�R�޶g���V,
�O������ba���w��D�Ƙ�2����I�����*�

����������$N�
��Rs�� D|C����-��yn<5�\�K��@3F�f��7�e�I�|ݨD�g5��i��v0�8Z�M�2}@LL
����RQ�����OH�-��p9�|�z���=��qr�g�[%�p��O�DJK=�^��Z���2�gJX�܃�U��
�.�ջm[��S��Tƽ���W5�-�݄̭�QK�(��'Ŗ���ķ����iA�g
 �$��84�s����:�ppp�����O�I�a�> �<
JN� :?��j��j�W��ɘ��6Q�˕?��7$�Iky���Oα���*OK-�vs�/F~�n�L]Ҽ2�38,mU!wX�V�ǳ4A�q�R6\��d0���I��'�ΨNBb���.��SY�*h�2$����~���a��jsܧ%,>h����_!}��:�5����A�C�NMn}O��&-&�ڤVA��p�~]��ث��H�ec�P������7�I��*�!� �@>%bP6�9ۗ�R��Z��@f����I���C���CUT{g��c7,-z�G��))cWR.��/�����W��c���4��Q��/�+R��{_d�0����qt̍`F����n�0w2��h�RQ8]��p�����������J����������v����V.�j����hFF��d�b/\ ��-����z�9�s�6Y��mt��vNTT�4�ӊi���݆��!O��vO�,����'e�]�%11_��I���*���������Ϙ�F�3&�%\y��գ�9\�X�&L� _�D�dՅ]D���qֽ �<�;�d��D��r=�v�B:�cGF�T�|��4_��8�4�,\�br��4����Y�E�d/�UC'��G�M�+I�I�I�hu`��&9i૏?�S<�?��B��N��T�ײ�V����<��~�~���9���u�V����$A���o��=���%�7�����_��@��� d%�LF�q����y��px	��ɪ�!�ѐ�G��w�?SA�
�����HH�����H�RLMOk�8܇?�WA��E������GD0sp0��gǂ�6.��PB`/,�dP=�M�ɠ�l_�M�/����u7r���0U����R�Y��$��C�+�����B_�@����� [o^	W�[u��6�|U�����k�{*ZzUv؃��x�]�[�GC��nʽy\��YY��|}��V;���"u��:�YG�J�cji���AX{C��]	8:`p��hm����f�j��r��[-�'}|(��n�&��0.���l9���^�FO��;3B}�b1��Zo�*j9��uqv�86Rr;ڗ!��7:��M$�=��۵�Z[e��W�J��x�C�������O��G��f�~����U��>X�"# y�o�=�O�'�b4�Eq�C�f7���^s21���`�*�8��h�S$��4뉭o��n'�
uv�x��Odz�����Tx{�~���6�xjhpY�:�8�uIlC�╿�	Z���$���@v ���MWu�0�P��b"���;~��v�tN��鳈v'Q�9#g��Y���+�����'�^'ly�klM�����Z�m�����WV~}��U��ة]=�q��DwF�]������D<�q��Ūw�f�&ox:���H��4v|T�aU�
L9@�H%E�,�fd����au�p�
z��R����0��1��31g�-Pv9�4�ת�������oMQ�x&���6�Bh�yy�񧟐I
���j����4l��։�F��Z�/�V|)5�ˆ��T�.�����>wD��Nl;�i���'荖��f�@LmO-�N���#T�J������eSw�`c��ߵ�Y���#5�c��"���7�O�4��}~�s���h�
�{�vC|�2wEu��v����r�㒲#����ѯ���P�.���yG�vr�i���ƺ�N?���֣N-n���I�z�#�j���|�(e�ٜ�6�J�6�=R�[�Wv�?o=�\0l�7ɩ��:���"`��zV�Ɯe����	��
�G���8WdǏ�eT�]��S�z9��]٩��0�Ē?���z�)|��;�I��M1�9�յ!3�`��,��x��'H
 �R�eE\��:(��l\�l�]r���옉�R�Ȕ������юWg0���1�ɜ���R<�X���v��c�;uk?ҏ��[�HN�����U�����P�WD�FL��?ٙŔ��&�Z3�$޳0��ށ�R:�
j�˹4�KCP#Jb$�����L��1�C�i���J�oS����,�9W�~��
��Z��o��Jl{⮂U��^CP� mzNV���Z=���7b��32���*_5#��.|��W"��2!d ݾ9k~�Ӹ1�;������uk�hW:kT��R�-�bV���(R����ѓ[Z��EG�r�n�2��t�1��6]ي^����PEɆI��M����*����}t����y����	��r�O�����8��Yߜ��O*Jqv�:/M> ����k-�W���M�Qv�kYI��O)���>"�̫:��L�
��}2Ha��4�X\^c=����B��/�G (&6&�͏�L86��*!��TF�삜�?��'�� �/A��|��C<]UPX���ݗ����m8zv�a2�؛tx���w��)&r�y{���܎��x�-�e�����_�I���W�x�\@�����:	zvvv>~����`8���a&P����===/Q_T�_*l�v>����Q��%��;3���n�C�CD�w˩h<+m�����%m�9����hpƀ������[��j;3��G_cϲ��������3:�ERo�/;��w����`c\ik'pC�����!K�L�	�Zp��y��eWJmNy�bXp�)�*��<���%�0�kɖ�I;FO���h :՟Z��ߙḸ�@�>��{z�^��hq)���p@��^y0.	��v��ڰ��m��":��50A�韙��Nj?I���RJ�r��Q�<g�o��1�}����jw�gk��(��܎���{Y�?��joDK��j�[	����s���qK��!����pK�J�J`�Ρ$u�FSY��&�&C�Z��GJ�#9�[��(�����7W9˙��%�S�Z	S
�?<��I��}x�pmg�I��=�͋,��D���K�yB�	NH ��L�zY�|=��H�r�Li�.��WoG���o֝y��.��>�������G�aE�*\`.`|-Fp6-ur6��#��D
333�tr��]�fML�"���Q{�G�������	YY�xmͫ�C##]��Q�ko����^9���zs2���f�쪣��L��>8�A�Co"��D)Q�ޘ���!�ڷ� +�d��\y<wI��ı��6�<�"�7Xg�0�Q�2)�)p�,w��/��YRNR���W��\��$��5���G#���1��r�7��NL�,��@�1){�嬅`:�����>�gYFYY�*��~��GK�(�ֳg#�wF���FWT$LdT�C�i��TGO��pO k+�@�v����-ߏ����54�@͔9��?�i��h8_I�>}3@p�=������!��CŖz���G�_疿�#�q�Z����)o8V�cA`~��_�Y�-,h��??��]���;�������2�oB��ctt4�?\$�h��5�A񱰲�oɝ�]u^-P���-�^������66dG![�5���nc�y�L�)����C���TJ ?�og!���V����Y~V��@$_�ɑ<�#�T"��R�i�n�͘�9ĝ'�z�1��Tl�qʻ����$<ߒ�
�Խ�z!����%���&7��$���������������)c�.(3�?1��
�;�}(���)���w�ȇ����H���\����x��uT~��B�Y˓_��M�>�n��/�����9=K��I��Ye8�� ?�k�p�;'��x�t�Q|Kr{=x�����&.�� H�yeeq�;�B�VF�����6��,�;|��{���i���*� ���TEAj��?������T�inE�_�K��5H�Q�����w��3s�3�Z��[1����J����.�� f�݋}�����M�"�<��@���R~��L@N�'4ڍ_Z�r���b��//���Q�w�����궣�C���2�W�^þ�3XCm���cOtt�ϽsT�P|�x�f�9 �.�I���\��/p��abIb<��̫�If��֣���|���d���������'��bٷ������f}��h�\�L��� �'/�(B�� �5�YR���]����=�S�B�9�h�N��4^��F���581D��^a�7�/V�@�F�@�{C�wL�Z(�̻rs'h�zg�Q�f���g�6���t99]����
D/d%��J)A��E�~j8v��x30Oӽ'��4���?O��<ܺ�c��vߍ�p��O������>7p�s`��3%�m\��9�U���s�J���B�4�!�]����n��f9��p9�8���ogDj�ne����JƋ/��M�..<�E�edd�L���'K`��$A �3�G�ffzo�2ʈj����ﻅ�Ay+�	r; '��	� .��@ˡE��~g�P���IG>L�0�B�N�rI�+�����P��x�{cZ�0\튬{�ʟ玗GD�	�L٥��4a��9X����>�-�{�!*:?��̓��믒g��2�'��P]��:����o�r�^i	��}s{ž�r���"�Y��h�juM�N��������+�qp�/;�!N�����ف����J[�z�]��������%N�To�D���_�C �����[�u��o9���.̜���{��3`��[_߽�]-��@]6�7T�����"�6.��Zv3m�t*�	S��_�y����e��׷�;�q&pR,����
 ��gx�*c��{�xŏ�\]0u�[t�8�WhWj'�C*�Z�ĵt����l#|�)�`d���v�t��F���:&�:���cE�`�q�d�c(� �>���EJ�
ݬ�Ь&�ϳ��/�m�!#'W�E��؏U��� Ӻ����*����ՑuT�r<�wmDU����8��ٲܖ}��J0�N������zU���=�a�����B�cBO��ѯ4��k��*%�X�D$�-GO;��lِ���a�w؛2O����ُ��V�s� �rZ)�U����jZNff�4���L_�4C�!����PÂ����o�Ҳ���:>52oq��ˈU��f&�s�tq1��NM���v<���j,Ur3*��a�׾����hRlm����(�N5������~�Q�VX�ղzv�	'�$��En5�����&�!��)�)VA��U��g�]Q�^���PN�u��>�r�}u�9��&�?�m���4AOqΰ.�;�ѝ��^��/�Uݼ��TA��>f������[Y�5]����)����m����)M�)�i+�]���¹��Z�u]��n��ͣ`k@�\�Vdí�����{-�k!-�y���x�2s즛��{mO�8�.�{Ng/G�����i9M���[�`j�Z��Qy��s6�Y^��:6��7�=&����S�/���e#XB����.����O�d)%m]t&"��ya��Cg�Ax�]'jGM�\^��	w�T\O��Me��`�͜T��k�n9Ӻ*p��"��H$A�x�GEf"�$�%�Mkn����s��x��h�D��8A������o7,������h��Q�Z�z�'w�vG �	��
���MzuVA�DM�W���H<���v�Y�k�����zB�OX���4~�e���Ҭ�QJ�~Y���/��6GLJI;�)��1nv3�+�$%�T�Ñ��+**2qr�7������V��������Ұ���h�]V��{���#��>R"��*�ؘҴO�[^z�l-͸!Jt������u�d����q�ɧ,B6�ga����-R!��O�ֲc~5N�?
z���ǟ��'�l�k�"(�`�DL��t��oQ9��,v�����2��i�Mp�h��nRO�WF�o�>�e��� V*�ga��b�P����ډ��R�����������(٩�S�
]�aX$Q�ֺ����8�մq�M�Šf����+Q�lx�p��M�S��u�|�*�t7��DU���ۘx.�%z0�.:.��Γ����lN�E�߭�陋�qa�z�Rđ�E��A�$`�>����,��B��4���̌�V��̈����mzvUUb��J��IX���\0l�Q��񫪆[it]�k����g{�cE�w��� Oj���J.��M�GJJ*��.�Wf,n%	�c��nud�eS���4��O����wiqvR-m��$�0��\_��0zy��`E������Ȃ�p��	�-`U���N2�/�j�tِ���	�3_#p~p���}���A:;�`����A'X��^��ӏǎ��(~]*0����Ԙ԰ށ��F�<��#ܳ�G��w#*n.w�-��SR8tnx�e����Tz{��D����U���r�}���b8�E��@G<$�9���22>��N�����i�:�:�ظ0
(<�\/�������g�bnptc���u�3U��Dܾ��Ŷ:W�|�!\]#x]��{6F��U���0j'#�1&��!����$�`���*�=���Ǹ����ۧ����=588}�ݘ&���`|����2���q��Z�!\3�NW�2c�3r���v�����L����\h�dG�;����SJ3>�פ��!��Lx��gH��E�*�����&�+�ǁ��XrQ��l�&O�CR�a�������LN���ʽ�4 .k{���u��wB��J>"�C�y�A>��B���)�JٽL들4L�V��Q�]���d5�{�`�53���!*��D&���7*~�������[=\�����N��q�KA����O��1�+˄�s����	�E<ùP7�bz���z�~YB6&�+����/�����~
�����g]b|%>8��FY��w|�!Y������t,rQ�(���#~N��Zڽ��=��L�{�Mu����~�{Y]Y���G��4T�N��8��jhC��dl7�w ����K&ƌL����֑AU�&���%�y_ s�m��\�P���΁ԝ_q���,�Q���i��=�����,xXW��H���g�$LKGpJ�Π<˙�����)�̣t��l��d��Srk�^&���4����Y���hKfc]r�ם-��P���=X�k�1sxdD�L�(gA>9k񙺳C�A�Uz�&v��t��n��%�7@��&�H�4�<�������'�:�l�wϢ<��� )#�?-��Ÿ[����oj�D@B�*�O���]������S�,xR-��[J����F�����~LʰI���vA�h�����U�Lܘ�}-�`k�,�����E{N]���I2O})A~m%LH���w��KN-]�󏆁N����S /^�6K���W?33�3vz�^����4���yJ��o���{�{�n�%0,s�i�q��N��(E�A �P���Y����w�fqSK��o���y�������O_^:�`��)�����і�9v�`�ez���/Or�>Q17�hJ/�q��ɢ4I���l�DUh�0���'zT�V��述�:��/�
$�)�f�6i���t?2��6��)S���R��VeX�)~��䭆v,[*I���E�P4��,�d�\��6����t�]�r��޼��A����M��lY�ؘ��jp�(n��m��L�o�;�����"*sP��0�0�4iZU�K������o�>q��n{�S�gG(~����l�_��򋛦�nܒ���8���v���}Vɓ�,rڜ��M �|˙���<ob�I�Ui7���vP]�Z�44`�wvd'�;�/��I�P_zݧ��L���t�
k�\L3f\����<����f)�O4������ntd����5�ԲLE;*Jed�8'�6�puP˭t�7���W�t�8��9d��E��
y�ڎY���6�8	8L�*)�Ö)��f=G/됧Q����5�c�鯃x�%p:K!�����_b|zҽ��g�ۥ���GSƌ��q�0w���݆#ڈ�tϢ�YG��=X��8Kva�,rބ�E�^X����~���n��Ә��@�M2�|���H�r��ھ��c�f���?�Q S�"�z��R2��޲_�����B�{waB2�Y�4-��}��X���֠C�-r�x��;:V�3>��>Yw������#}$��$�5b����K/���T7͜']c��X|��? ����i�554�U�JT�&�d����į�~�q3Ӹj'�B��o"�q:F���t.j!�����AD�X
��X��;����5�\��9�t�=�;�Nr��::j��b�6�sdZ籀� d��&�;��	����a)w�d~��dW����1PS�9*�� \��D
 ���s��xL��u��C���G�b�ZS��ߌi��y�}x�(�dc��eDMf܅�n:�� ������M@�����D���K]�fi�>����zF9��vפ�B^�=�:�����2cWl�3H�{�+V��E�$�_2��r^�$D�&��!��x��?�nc\���O�n���њ�yg��DS���:̓F��ǝ'�x�AJpx�=�_�{2Gr��ͺ�:U�g�S�F�Jh�j�(�ꖼ-|Wd��"�� ����Cu U:o���҅��?b�m�����0���e�4n��n���k�Ц�Ԧ�^�&Zң���LY����ʻ�:�Rz�P"6����\���f��*�l��}ɥ}��!뼖�8�nSI�mK�� 1���z�e\_�nM�ͭ�z�S�ٳ)�pHi��=��J�3w�~Ti���3���w�w���C�:F*<_�V膆ʡgޤpJ)/ݖ�č�Nt��S�Jbba�:��K��}u�n;�E}���F:��jH!pooo��//��F���h�y٦)��	�zA�_��\g�	k��ᆤt�o��6]�����Wϳ�g�{=�J���nH�|�/-�<�Ĥo�y6�7��m��no��T}||:���H;�3�e�R���߆�H�2�~ ][��1�RW�{��͍�%�BG��Ӂ���eL�(�,�ihW��$��B�sfj,�x��q�}��S��bJ~V.5F!�݃�s���h0�L�bjz�:�]>O��:�<!��;��7�V�e�ۯ�
��aiUP��y���R"[�͊2�sH��!#|R����0"Fn�#�-Q�wk))�c��緤	��q~��N;�Jt������4�:e�x����{��Fb$��t��1liI�VmY�!y��baa	l�AV;�u=���O'�X���V�,��l�'N�C���M�A��lE��7��?�#N~�{�
�A�m����b������9!��W��G5�z�H��W8_��m ��{z���bw��_ˣ]��`6p7ގ[Hw�To�]��R�CF&ҁ��U��_Ƥ����aT�v��/�Z�ॷ>�'���?MnY��G���M���{yB�U�;��vp���,7�v-�u�I�e��aw��n��_.�� �,�p<�������
9�P���mr��h���..�G a55�XZ�Ƣ��ʘ�\G�/FpNTzqF���Xj?�z����QF�;��Sj5H�{�N�����sa��f�y����Jr��=��o�^��jƦ��Ww�sc&{��*����0���E�<H24V�_���oe\k�#�5{�z���s�@����pʼ�#�[�����8�>g��2�[c�.��������[���3� ��k5��b����tbH�*Ɣ�U�����_%33��&ʴIQ���6+��2覫�B�<&����0{QQrޤՒ��e���2֦�v[�u2oQ�E�X�;�?}�?�L7Q�#��p��v��p�w`&M�� #@ܗ���)١8�<
'���EA���zwkS3��-�l��MW���V�\3%C�,R ��v�����k�k��x�����C$�ط�|^�aim��)��@��k��U�y�����f���l�h��a��6��w��c����Y��Ŏ���d���Ҵ�����i��D�"�>��&�yL���-�Ymp��vR��L4��ᛂ�\��c�3:��������+K�c ]�������f�|�[2 ��]T@�����h�@�Ͳ�5s�j���h�������ެ��q�f�J�'�U-W���ݳL^�J;���v�ma$|H�o���@ ��aʄ��=L��j�)TI��h��I);���jnE�"u�L��Q����_�u��
�v�%�4h�E����a�p�?="2��"���1�w��Q"8K�\Lk�62ĥ�w���:��q��sQQ�@BATVH�L�݋�7e�]��c-pʽ��4m 2�|*Y��%?���A2�v��Q9�Q��	qg�R����������q䡽B0�*M ����~�|]%/nHj�{lՑ�F�J]\gD4��@��/�y�/w�D�z�=���t������T#f&�m�@��d���'T�(��c	&�x�~�(*|���"DB �((j�W�eE�z���.�^��:`=ٙ�srr��%X@I	F��ͣ&7H��uw�?����\�>��*��YDٟW�~0�0S=T��� ��?f ��,��|_?)Y%�����b��l �K@�r���}��S+��J��_�ALz0� 0��F��ɷ`:4 ����qi���\] �x�3w�;�!-@W��=���%�Yϸ����Ԅl)��h��|7�:������7�%z#��n��B۝���A������!�+`(Yѫ=�*�����{9��i�e�Ab�K���o��oU_Xe}=������Z!���26.́��}�!���I�C�Y�:�N�$M�[R᮹�E}����qw�/_(��Kp}u�]O4���:�.�� ����/P��#3��������XM�u�����H4������]тs��F ���4��kߎ�ΆZ'8F�h����4Eb�K������'{]�
��q�k�jk8 �GW��Z�I=���|O�(b�FH+f�/��t��)	��"���Ƙ�ȕ��ːY?:]x��&�Ց�`9^��������+1X#ֈ�)�����y�Sj��c�/�@��'��V�YQn���޻4<މ��`ǁd�t��_!ԞXF��=�5@|*�(�p�.�L��Gw�]�1���"X��� [��) �cfg� 2Rd3�>��˯|�Z�6ͅ��S$�<�4tK���U��RwO�M�"T�e��� �G4���	�4/��*�&2��z��nFݷZR6X���cw���H�{���g���x2&KH�6�ř :[4n�0(j��.%�$$��QT?���z �{�R��`H����ē�=��Mco��>�y���6K��ᩁ���,��*)������Out�M�`Z9��xT�M��C����"�!�n��z���CHo�+́�K��?-R�t��S$���FO����M<]�=h�gqlM�'%�	@g%}|�C�lZ�[�PvJ��+@���������*+�(^H��WN��V%���n�}����}����Ms�9
���?lM�NT�&�8خ���.No5ʡ^k!���MڬK:����皣f �i�;�?��e�����G�'ZU][ (1N�D����Y������܏���K�����Z��	���z<�|/�	�B�ۜ�t��HoB��=4���� �B�'�p�,r�O@ �7OC@)������D/a�nD	YEy_�3�MU��˥�;�,�	��5�d�&�^�m�[泴0�j����Ɓ�d,�]N�Y�!d)y�)����zs�����ʊ�$V������`��/�:pt�f�srɥr��*|@���.�hii��K���Kp�g�?�y&93���� p�.����e�+��/�u�䔵��4���ʢ���l��%OE�ϼE;�)۠�; �P�G=����j�y膶�/�n3��uH����P��G+uL��]��			�GC�I�-�F_66X�.�W�l�_'���Ɉ���O�@\��,[\qߙ���3��ơ�sE�o�I�#x5��i����XԐ>�CU[X���;��5�
��O�?�:ޫ�$��`@��Y�|G�u�|���D( ��WG Z5�U�5���ku��>� ����4�A ر�9�{/�&�����#_�|��YA���Mw�r�o�wjЮ+���N����M�H�?�3����܅ќ���\~�+�f���b�j���;7�.�.[����� ��\d�ם��G�K��ԏ�����;�,���u�0��v5:�W�pbW멣���͏l@��c���N�]�f�27�ـ�h���l�U��s4�r�� ʨ�it�l����HԢ��)��.S�d�y�q�q~^"%5uȫ+��`��W�P�瀔6���\��M�}��x�׶晌�O�σ|� T7Hrk�1����B�~J��GD��FkF\�滳>��2��s���IG��L2���]�?��$�_���S-�\^C۞`� ����'brmy���@i���i!
μ=�,�p��W|wӄ��Ao�V~�K' A��_�޽��C�ô@�z a�@Y���>�5Ur��K]�ëBZ������� [e�%8�a����|�w�6�F�?_���#3� �t�f��QN��I=������<B�쎣���_�;[|o �8�4��H������?��݊�R_�4�Ê���gYz�Ԇ � 2%%�f[���e��c�U�6�+SD�*�K0J���kE�Dt�^�sv�����KA������߼�h�G
��蚵:U��P��蔶2j�S7�o�N| M(�1UM#�E��a:�����s7����r/�޾{�O��0��b 7? j�+z�����n���Qިר!Mٿ��@����}Y<}�`�������G ���Pŗ���%�!�w'\��ڵ'^�L߸!�Ď���U�+tnwץ�ރ<�}��W3k�:�DȢ��m�i�}�H�݅��!�S��� bz��/H]]v�eH2t�K%����svî�Of������[ ӮrO%������9�J:<�W+����d֣,�̔���%�}������k�������q�2�7_c���Q.F�  ���<Bq�n�9��|������9Y#
6���A�?z"9/:-���H�l�?�=���]�_�:����/��q�ht��[��5Q]QYy\��~�;��e�b��[��y�gd4^���T~��� `����ǱL��qF�w��2oWNGO���|t-��ZwJnT܆�e�2����ڕ�*!]wc�e��l@(zK�/܆�,������[��W��w�z<�G��6!�C'_i0$�8ѩ�w�f7�tq�yG'%�Bw� Qtf��%&>_��`��_v�4�uv���Uۋ ��E"U��YUP��(
ׄta7�Y���J�Ц����zw�L����W>�%��I#�j���⦖~����4��]�u�WG�E�B3� +��̶p�V�j��wG�_���) ��;>�7��;�&O�����I�_"�3��жzx<��&H�0�v��������q����]�,ж��l��{cH\�6	��X��k<��R��ı�?RO���R�s5�K�}.���%�M�k��wƦ��w���,��e����n��Q���z�3��B�T�Xm\%l����o���G��ă�����K^�ou�͗{B<��I����8�U�b�_W�LV����m�'~"��iP����կOKzs7�"����sf�K%���X~���`�WH�H$�+�۽��A����Q�r�j�����Y���.e�P-M�g$��$���+����F�yzߔ��& ��v��Si/m'�\"a�ubz�a��o98s0\h��\zz���^�f��p`F�}���tK��_w��4������ڲ��Z4��&���ة����~��9pN�驲�!���Q&<�	��b����pX�p�������a0(<���Ck
�Ơ��Ň��ǓBw��v��{��+xw-i'�_B
�Դ ���hʆۛ�wV��>���'z&�H)w7e��,���������L�|A��G�!�gg�!84<<�?+���,��hpEU������.�0�g�w�ȳ��nS.��ɸ��c�ļ�~�C&Їӝ�Wk�����&=`A�8��ӃV1�����{�l�����?�E3��G�o�ˡ�|��;^�#�����
��W�������ۋ�7�rw)$���̻�<삯z�^���'KFF��=}Ԣ��@�ѽ{�t�{�����Nvm�^���W�%���w���Sji�3܅��:_�Yd�������⻩���ƾ߬�6\�x]mDpr�I����@�����1kr�賄7�<���z�~�`�H���^�!F����g�B��m�spG��KC�<�\���h������\���s~���$�2���삇��/��2�����OG�ѳ��17�>��툢�Lw�����x(���O+E({B�lY'��C$�e�le��X�$K�Ad_BF����]H�=&cٷ��w����<������os��u�y�����:=������A~B����jQ�Ã'�?|1�X���Ў��}זN�䖄6���a�L��WGj�	/�;Y+dr6�WeRP���2��U�Y�����������w���o	��6q��;��	0�ԝqO��)��r��|�W�����7��NR�,E/Ɖ�H$	�0aҷ���=?2N��z����W4	�\u�.$�YY�h6��h��H�k|J����iҎI�XM��?�L�eC��71E�ſ����P�9��CU����ۀ y���d��'o�l�_z+,֧�3����0�B�M1�SN�}�I�;����=���П�z����������xP�&����Iokv�g%y�D �''pdk�߮��O=S�G����X&;a��yN��=�D@�C�=A��.M5�!�6���(��%��Ы�@p��ü�z.���\9�(Ϸc23���o ?�,�Eag��G5H� LVVv<�&�)�}T(Կ���A�f�:���]��[�ܦ���y��k`��P�|�_ŹU`z��p��Aڥ,�7���b'�#䗛�������������:�P��N����� E�)�+s�Շ��tC/&ĝV���=�Q���O���L���LpsB>2�\\��mlƂ�ޥX�#�c����?HG-�׸�7�FQa �5�5�1�EIb7	�n ����(��jn��+��y����z�5��;W�����g��y��/�� v����>sS&K�j���F�߯"��a�E?����d������4}��8Z,��E��ӧ~��i�P��?X�SS�фrʠ��a纲d���˕|�X�g�	�>�X�-I"�2�9� )��b&�3V�	d�w��Ɏ��"\�p񯱈�ÆqT�j����`y�ms�_�����|�h}O9�Q��o�M�C���"�ӊ�	m�f��/sS2h�N����?�-�I)��#��v�������|Ҕ��������@�7~�`\���sD�|e˥.K%��|W@䞴�"��D�4 j��i�Y.D��}ż�I��V�QtL��ўm��Q��Ϟrw�L�~r�����д��ۆ��:c�4h� ��;���gl�o	��1b9� S�^�z�h ,r�9�Z2����[DS�lU�U����7=��؍��oB9����w�}f��� ;).vN�DA0O�AQ7��+#m4M�e�#�O8�Gj���$��S+��'MLY񲷃��B���0y�����X[It��qH�^������?��v�l�l|��N�B�nwԭ6���Eee���U���M(SϽN-�Qo`�f��R�mx�?�%"�f�A�^�u*��3M�VssZ�w)	 ='H��/����~ ��͔�4Ҙ���i��a�= A��������:'�zR2#/c'�4�L�W@��Yy��V��5�8T������\�[�����u��z.�z�߭�d���7��'�sk{8�v%mHx�V�E ƅ�kK;28穟�,E���j?��	��*�[��'p6/XK�H�F���sJ�7����>zы�@�ؽ���k�j��L�{b1�����$����]]MnNk�ȿgב�~?M���n5��.�A�c�>�e�Ű�y9�&�:z("��e =��iV��q9_���:kOĨ�i�}�����Ѽ��9I��Ӫ9e��.Q����L�����.���g��f���X�cB�8���$}�n�"?��.�B�H�6��|�i2b.'Eωx��,�n1e�Mʻ��a�1�_�<�?�.E��x����8���Q��F�ڂW%5���Xox����~���i2���(;bc ��k���H�4��(��eB�͈��0��+�E9���=}:��6u|p��cd$�O�����k��$v#s�y��/�Y6�� M�/2�ӧ�R!�Ƞ�ҭ#��%�s2�3��m�.k��Ei�!+Lsb��3 )�I`���t�n��J����##�&�����;�
��d��q �gs�)YN�(�2����1�t+�	�m1��]22���y}�M�2ukw]t�|�&ٛ���)L1U��V�M�5V�e�e�v�u2�dԓnʃ�Դl�cv�����}�`�'�����a(q|��iR�x�ђ^䁖�XtS�V�J ��￨����"�;�.��$���P��v7>�VVa�;ޅ;��	��HU��I�{�[�)i6��)؆�:#ny7?N�Є�"�!/>�Ԥyc/��k�˩��t��Q�o��s?(��ݭ�ޡ�Co��aI W-��]�P��Y1���p��]���3Y��ʫ�}�(�����0����`O.d�ߨn/)�ɟ��&�m�Q`�y&Ho��l�MɯRŢ'�zxTu�.�"o%�8��.W8�n���W�k�[�x������D-쯆|Au[�l���RO̥���~[���V��œ���kqjӭq�����ǯﴈ�/R���z8|��L�v�L2{YS���PhM1Ϋ*R��S���h� �!���9�G����aD-#��))I�߉����|}���S��aL����#�i���	���p�v�M���wۢa�˻@�Wy
�H�4
�D���q�� ?Zˏ.�3�W\=T4��@�h�����Q�O�]iT�n�n���j�ܺ.�6��bys��L�R���W�:��!Gz�hx��0&v�����n+�L �5�/�4�"L|O��dq��N�P���w���|n&ӗ�����k�9:�H++k�p�K:��� �g^BTo��e�V������ ���x�8�(��f?۸ ��ށ�Ţ0li�IͽqW>C&���0���8�gR�'bx�NI�R]�r�ξu.�FA+++�D`�(�...�(}L���:.M� ` �:���E��n�C��f�qZ�����<گ�%g\��G%�w�:}�4�Ym�*xx��=���;������H���!�8i�H���v��cې}�z߈)m��L�@�^�C`��>�G?O{[]�'_^Y\���`0H !5�*2S&ZK��-__��v�F]��>gh�ډ��,��>ش��)��%GD���M���9G�fhe5����i$}�>������]��r�`��H-N��Tp�DX#���~�}�]D��'G-��)�ιb�{/m��׆�թdK7^��M�|�ў�`�uo�m�f`�����B��Rpǹq�T�e�[��R��G[Q�џ�P������y��4��NY��V�^�Rr���e�ʂ���Ga�z�s�.O��R�ȇ�i���);w���d�`���S�>��$0p܂Z-M��ˎ��w���u�S�GA�8mY�:��v;gs 2���ڞ�z�U�9���)�G-:^7������ ���6s������bClt+L�M�r�� 3�`�F���U��߻��kK����w�T��yP��L&���@*��O�Q�4^�\�P�5��q��s\��Nj��z�i�V�&��*4|���-~*h ���VJz<�8�ꘔ�F��W��-�K�����W"�'��:�� �)�]L��n��J�Gi*�"H�J,�3bQ~�����y9�Q����#f���2��߮%≬��N>�#[�>/'I.�6慲S4
s��3��R�p�e/��2���u��/��u0..grmʞ:��D�����=Z��&W��pǧ_��!K��$m��^]~�ꏩ(,(� �7�w<0�;�c|��P��.�8zb��c�Do$碈/4p4qtıʹ�D��0��]�w��H�_��,#|��R΃2�����Elӻ��D����ϐa��el���I�F ��[�Q<ӛ�Mv���`��/qv�w{^7yë�(A̯�-�=x�T�R��׿���.��-�׷��s��H\|�|�!���c.�W���F/���.�(��]T8��MW
u^?K�y�?jw���helL"����^�<����ҟ&g�x.°Ҿ= A�Lm(T䇯\]UUBmm��ʂ��w��+�ʪ6 TI�s�%r�E�K*��Pa�-w��E�q�*!z��˝�X��vv$)^��S�6̢�آ��2v�SCq��UF�ar�{��_����L���� ٯ�㖰��fY��c�D�.1
���mwD��ӄ,<�v���?n��A��Ɛ]������ E���w�&��s^^f_������bч�Y�&j�1��p��Qu�� �g�bр?4�7G��n��cE��7���Ԑi�:f+7�{�l�����i̵��\��~s�dӨ�r���-�M�qK���F]��� �s�BSk�w�`�2�J�����(F��'��[j��xuX>�@N�zu<�f{�R�����>S�kL@P�ZN�upﵴ���H��,#�1d�ý���n\Iz�vc>�q��+u�j��@>��)8��Xkn�^b��|�:>�QK9�:�|��ģ�TW9��S��Y���gsJ]�F�z�t^%����X�x�9q�2�=�>5��bK'T��k;����!��p��ə��6�Þ�/��|�%  �������
��&���F�R����z��M��� �y�߅�OŖ�/�V=h|N1}�xq��`��(P�mT}�-�@%���Ey1x��P(�����!�*�|�4L��Xf�ȆB�[SO��$h'EGKK<��Ե�>�N.y�F���u�7�>Mv5QHO����_�Tݼe�J\�(��]����V	4�p���miy���٩�TW��/�o�h�n���Gדg��9���ѻ�#^ll\<�e\h @k7O���BîY,0ޗ��j�j��n�*U��k�����dB��\������J�8]�-twe�"�8�&dS\F��X\w��~[��q�3y�cucv>�P����-����h����;���9����ro�K^��q����`�Su�`�[v���#�Od�:+�4`���H��c#;)�g_�Z�%�'KX��了0����Ս�D \�r��%[I4�f��}��̥��K����s�o�r�D�]�nuz�0�	w�+��"��,�G^�u�D�$���[V���_؉`:��г�;[%C��]�����D�@�e��_aK�Q��]�'l�����|����\h@܀�׵�Ţ���`�P�xpԥk
W ���i�{���-Τ�d�C��ثr�EƅWb#���21����t��հqVD�,�	& \�����H��ȝ�Ѻ:jn�e�7u
h'x"4�Xd�W�U& �0�	�,��W�%n#5n\u�Y��*��q9������k��"
�{02E��l��
��r�i�����Z?����+�˿{FT�S���{��t���{l�N����il�jLy���β�݈������Gʹ�fх:���)T.�Qw�FԲG��'��:U$QȈ����/�F�j�n٠����'-�c˕2.�+��z�lŝ9&��#���?[l��F+	����2�[	��P��"Nm�L��]������w�%��HC�	myov�� pUd��s�����@�}�b�Ԫ�,�蹸�u\�4
�MT�#�ɦ]�����y���)KD%����-�9�t���B�:%'	6��/h�iϾ�ZK��N�4m��u���W�u߫��U^8��zY��kqf!�c�yb��5�1	%.+W5�[��)&"�[_�z:��%�S䫩�a�k����
H���۪�ˬS�zh3(;`��{�?�F3�=Պ��=af�<8{���&n&�6Q�`�9�}�6h��L>�����u�Jc��n��4�r�����"e6Ҏo��-,�	N0�Qm�9h�AC�f��^�6�/H�6s&+!8����`���>���B!�\]�Q�E��.�a��6�I�㙪^���/\�Ƿ|?��ܳ���p?�T��,�|�h�����tdv���8�iߐ��r��vol�`&�,��I�:�x{̚�Г��(�i�sP�?� 0�ߡi�Ѧ�cR�y��r�ˎ/�&:/^���ր\�ؾ���d�+�=ov�U}�p�S>�줟s��c ]�-#�7:EIv� ��r	M�LA�uY�m�����^���4�y���=Z�������j��N�m����L�3��o��'�1�%�����լ����&���~�'^IW�fbZP"���r�^�$���"�R�V�2Ӯ��vN��kih�+�,M�M���2�P�]�3���]M�Z���`����ȥx?(H� 97Z��P4 c�0X��PE؈�z��V�dj�M�ge�gQb�~J�+��e�K�d`]i��/�E�.޸r�a��;� �-��E�����K�f��yy�O����7,�t-�ĉ[b?��e�.���_X5m_SP��Ԍv]�cW��_T�gl�ܱӬ'Ki�V�H�!�q�%�����+��c�IRJ��M�K���w�|�!�]��\T_[+a퉷/�v���B ��)#�K�e�T'�H
^6��ETw�����rA�6�O�ǜ�X7R��6~A��M�9d�0d��!�iji���5L�v��e���ݾ%n���O���v��+{5="7��x6V�x<��,Vl[k"�T	�l!Eʄ�~�9��/ �}eSH9nw�[���N5�����)�`D��U���$�8:�=>����!�D<ҽ� ��,E�j8hO,����{�S��RC�-�sn2��ۄ��/ͭ�e��\Q5G�+Z>qvu��~p��rt�n9(��a��gk��:7n��� �ŭ6UN��aY1l��Z��sRx��#��F, mZ!��*+�q=]�ˢԩ�gxrs���3�ˎ�r���}�+vB�����¿�Ֆ�[�E1���4]q���鼼�{FF6�m�KR{KS�u�ŉS������U������V��������Z-�?c6��l��s1� �DOTc.�[1bbhn���N���M}���.t0]E*�/d�͛��{iZ�!����|�[iy +������D��>}H#�g�M��E�x���,��� ��oN�� gsS��,�޲�~�پn�|t�Դ�p�~���.sӞWȎ��L�A\��_��b'}���s�i�^ַ������}�ƒk�=�i��sHn���ֻC�pf"&8�d3Rx����c\�A�E��и"U�u�a���Ӈh����]�:Q��ىBq^3CF������t�y�$��|�z쑳���I��Y��2��?�8�����յ����*�w�*Qث9"�/�I���*
�k��|nO�jwK?[���]
�9�\���ėRO18g:@{�tW�e�k���MI~&�w���7���g OxL��W��Yg���&7��7G�z=W�:H��Kk�˻����O1 |�/-}�X*���9�9�O9l��W��=��m�V)C9�N��K\�Ȉ�M��s`�"Rn�#�!M�w���~��w���)��WS�69y�ː_2�W�6��M����M���_���Pd�s���ۭ�DB��5=�����Ï�:&�軍�I
�b�	��4��)����y�p���Z	��$�ǉ�vu�"?��I��]���E���E���]G��E��ej�)���D)��y�����*���_��=M�;����PK   e*X�$M�  Q     jsons/user_defined.json��]o�6����ۙ�I�.���-�$�
� JTJ��<�N��;��4%���;K�s�����|�v�E�\�O�ߺ:_��|���	��d��q�_�����Ky?��6]�ID�Cf�~�_�w����:�����v���HgY��t�j$HY��I��Ve,�8�[/[/6�ֽ:�tC���f��O��U$��;ط���򋧼��/��^���w+�Ҝ����|w�}߽�Xr����˶��n���S}��=�!��n𣧟�
�
��P�T`e����m���a�˗�J�����ϋi6�g�9vS��7p4g!\�<���c}����524�r��ˀ�E*�×�,_|�̟�� n^�*���(��`�8���P�I�|n���N
�7��I��a�\}�+�!O2Gq��t7�����P���Q߭]���0���k�����[������ڡ��I���4� ZUH4L#�K�X#5�ת9��D�#�	�~�ݤ��A�Jo&�i��r!�c�8�L�*Ki(�(��Z��7�	=E��we3Y��J�$^���F���hM�&�rIU� �J�R�5rMC�\#Tu�&c��,�ц��	�c8��E)��/(�ce!���82��!����o(��ί���w}w��oj˭��$�"�@F�`� کF6��g�%!�!WvU*���vsH,�iV\+���a���:Ra^.��/1��'��
|�����$L�4�B�`����$΢�c����SS5Z�a��am�R�_��QE�׎׶BZ�
	�pd��t�S+;��G࣊��d�I'���I�X1Q�SFv�~ O]p&s+ð�_�S�;��ה}�q��y�Ľ�$�9������*S�	�V����ɓ@lR>�>�PK
   e*X���H&  C�                  cirkitFile.jsonPK
   p��W�C��B	 )	 /             u&  images/3fdb3be5-a051-4eb4-84dd-e907e6f5f8a3.pngPK
   ꩈWQ�O�  N�  /             0 images/5c74bc75-11cc-4f27-b1b5-62f572483d6f.pngPK
   ���W��W��: �: /             W� images/5eb2d398-7f6d-40aa-a255-437b4468b1bb.pngPK
   r��W�ѿ�*� �� /             � images/73de3dbc-74d6-4bf3-b63d-33bae631b402.pngPK
   O��W��ܣ]a  �d  /             �� images/7cd0bce8-56da-40c7-a6ad-eff1f7eef46c.pngPK
   e*X�$M�  Q               �^	 jsons/user_defined.jsonPK      S  _b	   